// --------------------------------------------------------------------
// Copyright (c) 2023 by JLSemi Inc.
// --------------------------------------------------------------------
//
//                     JLSemi
//                     Shanghai, China
//                     Name : Zhiling Guo
//                     Email: zlguo@jlsemi.com
//
// --------------------------------------------------------------------
// --------------------------------------------------------------------
//  Revision History:1.0
//  Date          By            Revision    Change Description
//---------------------------------------------------------------------
//  2024-05-14    zlguo         1.0         pulse_handshake
// --------------------------------------------------------------------
// --------------------------------------------------------------------
module pulse_handshake
(
    input   wire                        clk_in,
    input   wire                        rstn_in,
    input   wire                        vld_in,

    input   wire                        clk_out,
    input   wire                        rstn_out,
    output  wire                        vld_out
);

assign
endmodule
