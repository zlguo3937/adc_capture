# Created by MC2 : Version 2012.02.00.d on 2024/05/10, 14:39:04

#*********************************************************************************************************************/
# Software       : TSMC MEMORY COMPILER tsn28hpcpd127spsram_2012.02.00.d.180a						*/
# Technology     : TSMC 28nm CMOS LOGIC High Performance Compact Mobile Computing Plus 1P10M HKMG CU_ELK 0.9V				*/
#  Memory Type    : TSMC 28nm High Performance Compact Mobile Computing Plus Single Port SRAM with d127 bit cell HVT periphery */
# Library Name   : ts1n28hpcphvtb32768x18m16sso (user specify : TS1N28HPCPHVTB32768X18M16SSO)				*/
# Library Version: 180a												*/
# Generated Time : 2024/05/10, 14:38:57										*/
#*********************************************************************************************************************/
#															*/
# STATEMENT OF USE													*/
#															*/
# This information contains confidential and proprietary information of TSMC.					*/
# No part of this information may be reproduced, transmitted, transcribed,						*/
# stored in a retrieval system, or translated into any human or computer						*/
# language, in any form or by any means, electronic, mechanical, magnetic,						*/
# optical, chemical, manual, or otherwise, without the prior written permission					*/
# of TSMC. This information was prepared for informational purpose and is for					*/
# use by TSMC's customers only. TSMC reserves the right to make changes in the					*/
# information at any time and without notice.									*/
#															*/
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS1N28HPCPHVTB32768X18M16SSO
	CLASS BLOCK ;
	FOREIGN TS1N28HPCPHVTB32768X18M16SSO 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 654.735 BY 186.370 ;
	SYMMETRY X Y ;
	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 95.670 654.735 95.820 ;
			LAYER M1 ;
			RECT 654.555 95.670 654.735 95.820 ;
			LAYER M3 ;
			RECT 654.555 95.670 654.735 95.820 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[0]

	PIN A[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 85.810 654.735 85.960 ;
			LAYER M3 ;
			RECT 654.555 85.810 654.735 85.960 ;
			LAYER M2 ;
			RECT 654.555 85.810 654.735 85.960 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[10]

	PIN A[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 85.420 654.735 85.570 ;
			LAYER M2 ;
			RECT 654.555 85.420 654.735 85.570 ;
			LAYER M1 ;
			RECT 654.555 85.420 654.735 85.570 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[11]

	PIN A[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 98.110 654.735 98.260 ;
			LAYER M1 ;
			RECT 654.555 98.110 654.735 98.260 ;
			LAYER M3 ;
			RECT 654.555 98.110 654.735 98.260 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[12]

	PIN A[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 97.720 654.735 97.870 ;
			LAYER M1 ;
			RECT 654.555 97.720 654.735 97.870 ;
			LAYER M2 ;
			RECT 654.555 97.720 654.735 97.870 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[13]

	PIN A[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 96.060 654.735 96.210 ;
			LAYER M2 ;
			RECT 654.555 96.060 654.735 96.210 ;
			LAYER M3 ;
			RECT 654.555 96.060 654.735 96.210 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[14]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 94.010 654.735 94.160 ;
			LAYER M3 ;
			RECT 654.555 94.010 654.735 94.160 ;
			LAYER M2 ;
			RECT 654.555 94.010 654.735 94.160 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 93.620 654.735 93.770 ;
			LAYER M1 ;
			RECT 654.555 93.620 654.735 93.770 ;
			LAYER M2 ;
			RECT 654.555 93.620 654.735 93.770 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 83.760 654.735 83.910 ;
			LAYER M2 ;
			RECT 654.555 83.760 654.735 83.910 ;
			LAYER M3 ;
			RECT 654.555 83.760 654.735 83.910 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 89.520 654.735 89.670 ;
			LAYER M2 ;
			RECT 654.555 89.520 654.735 89.670 ;
			LAYER M1 ;
			RECT 654.555 89.520 654.735 89.670 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 87.860 654.735 88.010 ;
			LAYER M1 ;
			RECT 654.555 87.860 654.735 88.010 ;
			LAYER M3 ;
			RECT 654.555 87.860 654.735 88.010 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 87.470 654.735 87.620 ;
			LAYER M3 ;
			RECT 654.555 87.470 654.735 87.620 ;
			LAYER M1 ;
			RECT 654.555 87.470 654.735 87.620 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 91.960 654.735 92.110 ;
			LAYER M1 ;
			RECT 654.555 91.960 654.735 92.110 ;
			LAYER M3 ;
			RECT 654.555 91.960 654.735 92.110 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 91.570 654.735 91.720 ;
			LAYER M3 ;
			RECT 654.555 91.570 654.735 91.720 ;
			LAYER M2 ;
			RECT 654.555 91.570 654.735 91.720 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 89.910 654.735 90.060 ;
			LAYER M1 ;
			RECT 654.555 89.910 654.735 90.060 ;
			LAYER M3 ;
			RECT 654.555 89.910 654.735 90.060 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[9]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 99.770 654.735 99.920 ;
			LAYER M2 ;
			RECT 654.555 99.770 654.735 99.920 ;
			LAYER M1 ;
			RECT 654.555 99.770 654.735 99.920 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.115300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.228300 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.515900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.249900 LAYER M2 ;
		ANTENNAMAXAREACAR 10.191100 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.732500 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 11.091100 LAYER M3 ;
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 100.400 654.735 100.550 ;
			LAYER M3 ;
			RECT 654.555 100.400 654.735 100.550 ;
			LAYER M1 ;
			RECT 654.555 100.400 654.735 100.550 ;
		END
		ANTENNAGATEAREA 2.013900 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 3.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 5.372500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.331500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA1 ;
		ANTENNAGATEAREA 2.013900 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 2.694600 LAYER M2 ;
		ANTENNAMAXAREACAR 33.912400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.292500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.097200 LAYER VIA2 ;
		ANTENNAGATEAREA 2.013900 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 2.754400 LAYER M3 ;
		ANTENNAMAXAREACAR 35.107800 LAYER M3 ;
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 6.635 654.735 6.785 ;
			LAYER M1 ;
			RECT 654.555 6.635 654.735 6.785 ;
			LAYER M3 ;
			RECT 654.555 6.635 654.735 6.785 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[0]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 116.555 654.735 116.705 ;
			LAYER M2 ;
			RECT 654.555 116.555 654.735 116.705 ;
			LAYER M1 ;
			RECT 654.555 116.555 654.735 116.705 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 125.835 654.735 125.985 ;
			LAYER M1 ;
			RECT 654.555 125.835 654.735 125.985 ;
			LAYER M3 ;
			RECT 654.555 125.835 654.735 125.985 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 135.115 654.735 135.265 ;
			LAYER M1 ;
			RECT 654.555 135.115 654.735 135.265 ;
			LAYER M3 ;
			RECT 654.555 135.115 654.735 135.265 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 144.395 654.735 144.545 ;
			LAYER M1 ;
			RECT 654.555 144.395 654.735 144.545 ;
			LAYER M3 ;
			RECT 654.555 144.395 654.735 144.545 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 153.675 654.735 153.825 ;
			LAYER M3 ;
			RECT 654.555 153.675 654.735 153.825 ;
			LAYER M1 ;
			RECT 654.555 153.675 654.735 153.825 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 162.955 654.735 163.105 ;
			LAYER M1 ;
			RECT 654.555 162.955 654.735 163.105 ;
			LAYER M3 ;
			RECT 654.555 162.955 654.735 163.105 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 172.235 654.735 172.385 ;
			LAYER M3 ;
			RECT 654.555 172.235 654.735 172.385 ;
			LAYER M1 ;
			RECT 654.555 172.235 654.735 172.385 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 181.515 654.735 181.665 ;
			LAYER M1 ;
			RECT 654.555 181.515 654.735 181.665 ;
			LAYER M3 ;
			RECT 654.555 181.515 654.735 181.665 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[17]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 15.915 654.735 16.065 ;
			LAYER M1 ;
			RECT 654.555 15.915 654.735 16.065 ;
			LAYER M2 ;
			RECT 654.555 15.915 654.735 16.065 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 25.195 654.735 25.345 ;
			LAYER M1 ;
			RECT 654.555 25.195 654.735 25.345 ;
			LAYER M3 ;
			RECT 654.555 25.195 654.735 25.345 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 34.475 654.735 34.625 ;
			LAYER M1 ;
			RECT 654.555 34.475 654.735 34.625 ;
			LAYER M2 ;
			RECT 654.555 34.475 654.735 34.625 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 43.755 654.735 43.905 ;
			LAYER M3 ;
			RECT 654.555 43.755 654.735 43.905 ;
			LAYER M1 ;
			RECT 654.555 43.755 654.735 43.905 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 53.035 654.735 53.185 ;
			LAYER M2 ;
			RECT 654.555 53.035 654.735 53.185 ;
			LAYER M1 ;
			RECT 654.555 53.035 654.735 53.185 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 62.315 654.735 62.465 ;
			LAYER M2 ;
			RECT 654.555 62.315 654.735 62.465 ;
			LAYER M1 ;
			RECT 654.555 62.315 654.735 62.465 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 71.595 654.735 71.745 ;
			LAYER M3 ;
			RECT 654.555 71.595 654.735 71.745 ;
			LAYER M1 ;
			RECT 654.555 71.595 654.735 71.745 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 76.235 654.735 76.385 ;
			LAYER M3 ;
			RECT 654.555 76.235 654.735 76.385 ;
			LAYER M2 ;
			RECT 654.555 76.235 654.735 76.385 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 109.595 654.735 109.745 ;
			LAYER M2 ;
			RECT 654.555 109.595 654.735 109.745 ;
			LAYER M3 ;
			RECT 654.555 109.595 654.735 109.745 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[9]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 7.645 654.735 7.795 ;
			LAYER M1 ;
			RECT 654.555 7.645 654.735 7.795 ;
			LAYER M3 ;
			RECT 654.555 7.645 654.735 7.795 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[0]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 117.565 654.735 117.715 ;
			LAYER M3 ;
			RECT 654.555 117.565 654.735 117.715 ;
			LAYER M2 ;
			RECT 654.555 117.565 654.735 117.715 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 126.845 654.735 126.995 ;
			LAYER M2 ;
			RECT 654.555 126.845 654.735 126.995 ;
			LAYER M3 ;
			RECT 654.555 126.845 654.735 126.995 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 136.125 654.735 136.275 ;
			LAYER M3 ;
			RECT 654.555 136.125 654.735 136.275 ;
			LAYER M1 ;
			RECT 654.555 136.125 654.735 136.275 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 145.405 654.735 145.555 ;
			LAYER M2 ;
			RECT 654.555 145.405 654.735 145.555 ;
			LAYER M1 ;
			RECT 654.555 145.405 654.735 145.555 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 154.685 654.735 154.835 ;
			LAYER M2 ;
			RECT 654.555 154.685 654.735 154.835 ;
			LAYER M3 ;
			RECT 654.555 154.685 654.735 154.835 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 163.965 654.735 164.115 ;
			LAYER M2 ;
			RECT 654.555 163.965 654.735 164.115 ;
			LAYER M3 ;
			RECT 654.555 163.965 654.735 164.115 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 173.245 654.735 173.395 ;
			LAYER M2 ;
			RECT 654.555 173.245 654.735 173.395 ;
			LAYER M1 ;
			RECT 654.555 173.245 654.735 173.395 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 182.525 654.735 182.675 ;
			LAYER M1 ;
			RECT 654.555 182.525 654.735 182.675 ;
			LAYER M3 ;
			RECT 654.555 182.525 654.735 182.675 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[17]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 16.925 654.735 17.075 ;
			LAYER M1 ;
			RECT 654.555 16.925 654.735 17.075 ;
			LAYER M2 ;
			RECT 654.555 16.925 654.735 17.075 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 26.205 654.735 26.355 ;
			LAYER M3 ;
			RECT 654.555 26.205 654.735 26.355 ;
			LAYER M1 ;
			RECT 654.555 26.205 654.735 26.355 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 35.485 654.735 35.635 ;
			LAYER M3 ;
			RECT 654.555 35.485 654.735 35.635 ;
			LAYER M1 ;
			RECT 654.555 35.485 654.735 35.635 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 44.765 654.735 44.915 ;
			LAYER M3 ;
			RECT 654.555 44.765 654.735 44.915 ;
			LAYER M1 ;
			RECT 654.555 44.765 654.735 44.915 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 54.045 654.735 54.195 ;
			LAYER M1 ;
			RECT 654.555 54.045 654.735 54.195 ;
			LAYER M2 ;
			RECT 654.555 54.045 654.735 54.195 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 63.325 654.735 63.475 ;
			LAYER M2 ;
			RECT 654.555 63.325 654.735 63.475 ;
			LAYER M1 ;
			RECT 654.555 63.325 654.735 63.475 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 72.605 654.735 72.755 ;
			LAYER M3 ;
			RECT 654.555 72.605 654.735 72.755 ;
			LAYER M2 ;
			RECT 654.555 72.605 654.735 72.755 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 77.245 654.735 77.395 ;
			LAYER M3 ;
			RECT 654.555 77.245 654.735 77.395 ;
			LAYER M1 ;
			RECT 654.555 77.245 654.735 77.395 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 110.605 654.735 110.755 ;
			LAYER M2 ;
			RECT 654.555 110.605 654.735 110.755 ;
			LAYER M1 ;
			RECT 654.555 110.605 654.735 110.755 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[9]

	PIN SD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 81.145 654.735 81.295 ;
			LAYER M2 ;
			RECT 654.555 81.145 654.735 81.295 ;
			LAYER M3 ;
			RECT 654.555 81.145 654.735 81.295 ;
		END
		ANTENNAGATEAREA 0.051000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.839700 LAYER M1 ;
		ANTENNAMAXAREACAR 9.087800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.585600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.051000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.499900 LAYER M2 ;
		ANTENNAMAXAREACAR 48.990700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.878400 LAYER VIA2 ;
		ANTENNAGATEAREA 0.051000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.590600 LAYER M3 ;
		ANTENNAMAXAREACAR 48.990700 LAYER M3 ;
	END SD

	PIN SLP
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 81.860 654.735 82.010 ;
			LAYER M3 ;
			RECT 654.555 81.860 654.735 82.010 ;
			LAYER M1 ;
			RECT 654.555 81.860 654.735 82.010 ;
		END
		ANTENNAGATEAREA 0.027000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.172400 LAYER M1 ;
		ANTENNAMAXAREACAR 8.260000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.433300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.027000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.269000 LAYER M2 ;
		ANTENNAMAXAREACAR 48.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.027000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.564300 LAYER M3 ;
		ANTENNAMAXAREACAR 48.814800 LAYER M3 ;
	END SLP

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.000 4.875 654.345 5.205 ;
			LAYER M4 ;
			RECT 0.000 14.155 654.345 14.485 ;
			LAYER M4 ;
			RECT 0.000 23.435 654.345 23.765 ;
			LAYER M4 ;
			RECT 0.000 32.715 654.345 33.045 ;
			LAYER M4 ;
			RECT 0.000 41.995 654.345 42.325 ;
			LAYER M4 ;
			RECT 0.000 51.275 654.345 51.605 ;
			LAYER M4 ;
			RECT 0.000 60.555 654.345 60.885 ;
			LAYER M4 ;
			RECT 0.000 69.835 654.345 70.165 ;
			LAYER M4 ;
			RECT 0.000 79.115 654.735 79.445 ;
			LAYER M4 ;
			RECT 0.000 91.755 654.735 92.325 ;
			LAYER M4 ;
			RECT 0.000 92.455 654.735 93.025 ;
			LAYER M4 ;
			RECT 0.000 99.435 654.735 100.005 ;
			LAYER M4 ;
			RECT 0.000 105.515 654.735 105.845 ;
			LAYER M4 ;
			RECT 0.000 114.795 654.345 115.125 ;
			LAYER M4 ;
			RECT 0.000 124.075 654.345 124.405 ;
			LAYER M4 ;
			RECT 0.000 133.355 654.345 133.685 ;
			LAYER M4 ;
			RECT 0.000 142.635 654.345 142.965 ;
			LAYER M4 ;
			RECT 0.000 151.915 654.345 152.245 ;
			LAYER M4 ;
			RECT 0.000 161.195 654.345 161.525 ;
			LAYER M4 ;
			RECT 0.000 170.475 654.345 170.805 ;
			LAYER M4 ;
			RECT 0.000 179.755 654.345 180.085 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.000 6.285 654.345 6.665 ;
			LAYER M4 ;
			RECT 0.000 15.565 654.345 15.945 ;
			LAYER M4 ;
			RECT 0.000 24.845 654.345 25.225 ;
			LAYER M4 ;
			RECT 0.000 34.125 654.345 34.505 ;
			LAYER M4 ;
			RECT 0.000 43.405 654.345 43.785 ;
			LAYER M4 ;
			RECT 0.000 52.685 654.345 53.065 ;
			LAYER M4 ;
			RECT 0.000 61.965 654.345 62.345 ;
			LAYER M4 ;
			RECT 0.000 71.245 654.345 71.625 ;
			LAYER M4 ;
			RECT 0.000 80.525 654.735 80.905 ;
			LAYER M4 ;
			RECT 0.000 90.355 654.735 90.925 ;
			LAYER M4 ;
			RECT 0.000 91.055 654.735 91.625 ;
			LAYER M4 ;
			RECT 0.000 93.385 654.735 93.955 ;
			LAYER M4 ;
			RECT 0.000 106.925 654.735 107.305 ;
			LAYER M4 ;
			RECT 0.000 116.205 654.345 116.585 ;
			LAYER M4 ;
			RECT 0.000 125.485 654.345 125.865 ;
			LAYER M4 ;
			RECT 0.000 134.765 654.345 135.145 ;
			LAYER M4 ;
			RECT 0.000 144.045 654.345 144.425 ;
			LAYER M4 ;
			RECT 0.000 153.325 654.345 153.705 ;
			LAYER M4 ;
			RECT 0.000 162.605 654.345 162.985 ;
			LAYER M4 ;
			RECT 0.000 171.885 654.345 172.265 ;
			LAYER M4 ;
			RECT 0.000 181.165 654.345 181.545 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 83.370 654.735 83.520 ;
			LAYER M3 ;
			RECT 654.555 83.370 654.735 83.520 ;
			LAYER M1 ;
			RECT 654.555 83.370 654.735 83.520 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.445400 LAYER M2 ;
		ANTENNAMAXAREACAR 16.888300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 17.788300 LAYER M3 ;
	END WEB

	OBS
		# Promoted blockages
		LAYER M2 ;
		RECT 654.555 77.475 654.735 81.065 ;
		LAYER M3 ;
		RECT 654.555 71.825 654.735 72.525 ;
		LAYER VIA3 ;
		RECT 654.555 71.825 654.735 72.525 ;
		LAYER M1 ;
		RECT 654.555 71.805 654.735 72.545 ;
		LAYER M1 ;
		RECT 654.555 145.615 654.735 153.615 ;
		LAYER M3 ;
		RECT 654.555 145.635 654.735 153.595 ;
		LAYER VIA3 ;
		RECT 654.555 145.635 654.735 153.595 ;
		LAYER M2 ;
		RECT 654.555 145.635 654.735 153.595 ;
		LAYER VIA3 ;
		RECT 654.555 77.475 654.735 81.065 ;
		LAYER M3 ;
		RECT 654.555 77.475 654.735 81.065 ;
		LAYER M1 ;
		RECT 654.555 144.605 654.735 145.345 ;
		LAYER VIA3 ;
		RECT 654.555 81.375 654.735 81.780 ;
		LAYER M2 ;
		RECT 654.555 81.375 654.735 81.780 ;
		LAYER M3 ;
		RECT 654.555 81.375 654.735 81.780 ;
		LAYER M2 ;
		RECT 654.555 83.600 654.735 83.680 ;
		LAYER M3 ;
		RECT 654.555 83.600 654.735 83.680 ;
		LAYER VIA3 ;
		RECT 654.555 83.600 654.735 83.680 ;
		LAYER M1 ;
		RECT 654.555 83.580 654.735 83.700 ;
		LAYER M2 ;
		RECT 654.555 83.990 654.735 85.340 ;
		LAYER M3 ;
		RECT 654.555 83.990 654.735 85.340 ;
		LAYER VIA3 ;
		RECT 654.555 83.990 654.735 85.340 ;
		LAYER M2 ;
		RECT 654.555 86.040 654.735 87.390 ;
		LAYER M3 ;
		RECT 654.555 135.345 654.735 136.045 ;
		LAYER VIA3 ;
		RECT 654.555 135.345 654.735 136.045 ;
		LAYER M2 ;
		RECT 654.555 135.345 654.735 136.045 ;
		LAYER M1 ;
		RECT 654.555 82.070 654.735 83.310 ;
		LAYER VIA3 ;
		RECT 654.555 82.090 654.735 83.290 ;
		LAYER M1 ;
		RECT 654.555 83.970 654.735 85.360 ;
		LAYER M2 ;
		RECT 654.555 82.090 654.735 83.290 ;
		LAYER M3 ;
		RECT 654.555 82.090 654.735 83.290 ;
		LAYER M3 ;
		RECT 654.555 144.625 654.735 145.325 ;
		LAYER M2 ;
		RECT 654.555 144.625 654.735 145.325 ;
		LAYER VIA3 ;
		RECT 654.555 144.625 654.735 145.325 ;
		LAYER VIA3 ;
		RECT 654.555 136.355 654.735 144.315 ;
		LAYER M1 ;
		RECT 654.555 85.630 654.735 85.750 ;
		LAYER M3 ;
		RECT 654.555 85.650 654.735 85.730 ;
		LAYER M2 ;
		RECT 654.555 85.650 654.735 85.730 ;
		LAYER M1 ;
		RECT 654.555 86.020 654.735 87.410 ;
		LAYER VIA3 ;
		RECT 654.555 86.040 654.735 87.390 ;
		LAYER M3 ;
		RECT 654.555 86.040 654.735 87.390 ;
		LAYER M1 ;
		RECT 654.555 109.805 654.735 110.545 ;
		LAYER M1 ;
		RECT 654.555 116.765 654.735 117.505 ;
		LAYER M1 ;
		RECT 654.555 117.775 654.735 125.775 ;
		LAYER M2 ;
		RECT 654.555 127.075 654.735 135.035 ;
		LAYER M2 ;
		RECT 654.555 100.630 654.735 109.515 ;
		LAYER M1 ;
		RECT 654.555 100.610 654.735 109.535 ;
		LAYER M1 ;
		RECT 654.555 127.055 654.735 135.055 ;
		LAYER M3 ;
		RECT 654.555 54.275 654.735 62.235 ;
		LAYER M2 ;
		RECT 654.555 53.265 654.735 53.965 ;
		LAYER VIA3 ;
		RECT 654.555 53.265 654.735 53.965 ;
		LAYER M3 ;
		RECT 654.555 53.265 654.735 53.965 ;
		LAYER M1 ;
		RECT 654.555 62.525 654.735 63.265 ;
		LAYER M2 ;
		RECT 654.555 63.555 654.735 71.515 ;
		LAYER M3 ;
		RECT 654.555 43.985 654.735 44.685 ;
		LAYER M3 ;
		RECT 654.555 62.545 654.735 63.245 ;
		LAYER M3 ;
		RECT 654.555 63.555 654.735 71.515 ;
		LAYER VIA3 ;
		RECT 654.555 62.545 654.735 63.245 ;
		LAYER M2 ;
		RECT 654.555 62.545 654.735 63.245 ;
		LAYER M1 ;
		RECT 654.555 43.965 654.735 44.705 ;
		LAYER M1 ;
		RECT 654.555 35.695 654.735 43.695 ;
		LAYER M2 ;
		RECT 654.555 44.995 654.735 52.955 ;
		LAYER M3 ;
		RECT 654.555 44.995 654.735 52.955 ;
		LAYER M1 ;
		RECT 654.555 44.975 654.735 52.975 ;
		LAYER M2 ;
		RECT 654.555 43.985 654.735 44.685 ;
		LAYER VIA3 ;
		RECT 654.555 43.985 654.735 44.685 ;
		LAYER M1 ;
		RECT 654.555 25.405 654.735 26.145 ;
		LAYER M2 ;
		RECT 654.555 35.715 654.735 43.675 ;
		LAYER M3 ;
		RECT 654.555 35.715 654.735 43.675 ;
		LAYER VIA3 ;
		RECT 654.555 35.715 654.735 43.675 ;
		LAYER M2 ;
		RECT 654.555 54.275 654.735 62.235 ;
		LAYER VIA3 ;
		RECT 654.555 54.275 654.735 62.235 ;
		LAYER M1 ;
		RECT 654.555 53.245 654.735 53.985 ;
		LAYER M2 ;
		RECT 654.555 89.750 654.735 89.830 ;
		LAYER M1 ;
		RECT 654.555 89.730 654.735 89.850 ;
		LAYER M2 ;
		RECT 654.555 88.090 654.735 89.440 ;
		LAYER VIA3 ;
		RECT 654.555 88.090 654.735 89.440 ;
		LAYER M3 ;
		RECT 654.555 89.750 654.735 89.830 ;
		LAYER VIA3 ;
		RECT 654.555 89.750 654.735 89.830 ;
		LAYER M1 ;
		RECT 654.555 88.070 654.735 89.460 ;
		LAYER M2 ;
		RECT 654.555 87.700 654.735 87.780 ;
		LAYER M1 ;
		RECT 654.555 87.680 654.735 87.800 ;
		LAYER M3 ;
		RECT 654.555 88.090 654.735 89.440 ;
		LAYER VIA3 ;
		RECT 654.555 85.650 654.735 85.730 ;
		LAYER M3 ;
		RECT 654.555 109.825 654.735 110.525 ;
		LAYER VIA3 ;
		RECT 654.555 109.825 654.735 110.525 ;
		LAYER M2 ;
		RECT 654.555 109.825 654.735 110.525 ;
		LAYER M3 ;
		RECT 654.555 100.630 654.735 109.515 ;
		LAYER VIA3 ;
		RECT 654.555 100.630 654.735 109.515 ;
		LAYER M3 ;
		RECT 654.555 87.700 654.735 87.780 ;
		LAYER VIA3 ;
		RECT 654.555 87.700 654.735 87.780 ;
		LAYER M1 ;
		RECT 654.555 77.455 654.735 81.085 ;
		LAYER M1 ;
		RECT 654.555 81.355 654.735 81.800 ;
		LAYER M2 ;
		RECT 654.555 90.140 654.735 91.490 ;
		LAYER M2 ;
		RECT 654.555 92.190 654.735 93.540 ;
		LAYER M1 ;
		RECT 654.555 92.170 654.735 93.560 ;
		LAYER M1 ;
		RECT 654.555 91.780 654.735 91.900 ;
		LAYER M3 ;
		RECT 654.555 90.140 654.735 91.490 ;
		LAYER VIA3 ;
		RECT 654.555 90.140 654.735 91.490 ;
		LAYER VIA3 ;
		RECT 654.555 91.800 654.735 91.880 ;
		LAYER M2 ;
		RECT 654.555 91.800 654.735 91.880 ;
		LAYER M3 ;
		RECT 654.555 91.800 654.735 91.880 ;
		LAYER VIA3 ;
		RECT 654.555 92.190 654.735 93.540 ;
		LAYER M3 ;
		RECT 654.555 92.190 654.735 93.540 ;
		LAYER M1 ;
		RECT 654.555 93.830 654.735 93.950 ;
		LAYER M2 ;
		RECT 654.555 93.850 654.735 93.930 ;
		LAYER VIA3 ;
		RECT 654.555 93.850 654.735 93.930 ;
		LAYER M3 ;
		RECT 654.555 93.850 654.735 93.930 ;
		LAYER M2 ;
		RECT 654.555 34.705 654.735 35.405 ;
		LAYER M1 ;
		RECT 654.555 34.685 654.735 35.425 ;
		LAYER M3 ;
		RECT 654.555 26.435 654.735 34.395 ;
		LAYER M2 ;
		RECT 654.555 26.435 654.735 34.395 ;
		LAYER VIA3 ;
		RECT 654.555 44.995 654.735 52.955 ;
		LAYER M1 ;
		RECT 654.555 54.255 654.735 62.255 ;
		LAYER M2 ;
		RECT 654.555 25.425 654.735 26.125 ;
		LAYER M3 ;
		RECT 654.555 25.425 654.735 26.125 ;
		LAYER VIA3 ;
		RECT 654.555 25.425 654.735 26.125 ;
		LAYER M2 ;
		RECT 654.555 16.145 654.735 16.845 ;
		LAYER M1 ;
		RECT 654.555 16.125 654.735 16.865 ;
		LAYER M2 ;
		RECT 654.555 6.865 654.735 7.565 ;
		LAYER M3 ;
		RECT 654.555 6.865 654.735 7.565 ;
		LAYER M1 ;
		RECT 654.555 17.135 654.735 25.135 ;
		LAYER VIA3 ;
		RECT 654.555 17.155 654.735 25.115 ;
		LAYER M1 ;
		RECT 654.555 0.000 654.735 6.575 ;
		LAYER M2 ;
		RECT 654.555 0.000 654.735 6.555 ;
		LAYER M3 ;
		RECT 654.555 0.000 654.735 6.555 ;
		LAYER VIA3 ;
		RECT 654.555 0.000 654.735 6.555 ;
		LAYER VIA3 ;
		RECT 654.555 34.705 654.735 35.405 ;
		LAYER M3 ;
		RECT 654.555 34.705 654.735 35.405 ;
		LAYER VIA3 ;
		RECT 654.555 26.435 654.735 34.395 ;
		LAYER M1 ;
		RECT 654.555 26.415 654.735 34.415 ;
		LAYER M3 ;
		RECT 654.555 16.145 654.735 16.845 ;
		LAYER VIA3 ;
		RECT 654.555 16.145 654.735 16.845 ;
		LAYER VIA3 ;
		RECT 654.555 6.865 654.735 7.565 ;
		LAYER M3 ;
		RECT 654.555 95.900 654.735 95.980 ;
		LAYER VIA3 ;
		RECT 654.555 95.900 654.735 95.980 ;
		LAYER M1 ;
		RECT 654.555 94.220 654.735 95.610 ;
		LAYER M1 ;
		RECT 654.555 95.880 654.735 96.000 ;
		LAYER VIA3 ;
		RECT 654.555 94.240 654.735 95.590 ;
		LAYER M2 ;
		RECT 654.555 94.240 654.735 95.590 ;
		LAYER M3 ;
		RECT 654.555 94.240 654.735 95.590 ;
		LAYER M3 ;
		RECT 654.555 97.950 654.735 98.030 ;
		LAYER M2 ;
		RECT 654.555 97.950 654.735 98.030 ;
		LAYER VIA3 ;
		RECT 654.555 97.950 654.735 98.030 ;
		LAYER VIA3 ;
		RECT 654.555 96.290 654.735 97.640 ;
		LAYER VIA3 ;
		RECT 654.555 100.000 654.735 100.320 ;
		LAYER M1 ;
		RECT 654.555 99.980 654.735 100.340 ;
		LAYER M3 ;
		RECT 654.555 98.340 654.735 99.690 ;
		LAYER VIA3 ;
		RECT 654.555 98.340 654.735 99.690 ;
		LAYER M1 ;
		RECT 654.555 90.120 654.735 91.510 ;
		LAYER M3 ;
		RECT 654.555 100.000 654.735 100.320 ;
		LAYER M2 ;
		RECT 654.555 96.290 654.735 97.640 ;
		LAYER M3 ;
		RECT 654.555 96.290 654.735 97.640 ;
		LAYER M1 ;
		RECT 654.555 96.270 654.735 97.660 ;
		LAYER M2 ;
		RECT 654.555 95.900 654.735 95.980 ;
		LAYER M1 ;
		RECT 654.555 98.320 654.735 99.710 ;
		LAYER M2 ;
		RECT 654.555 98.340 654.735 99.690 ;
		LAYER M1 ;
		RECT 654.555 97.930 654.735 98.050 ;
		LAYER M2 ;
		RECT 654.555 100.000 654.735 100.320 ;
		LAYER M4 ;
		RECT 654.345 102.370 654.735 105.515 ;
		LAYER M1 ;
		RECT 654.555 110.815 654.735 116.495 ;
		LAYER M2 ;
		RECT 654.555 116.785 654.735 117.485 ;
		LAYER M3 ;
		RECT 654.555 116.785 654.735 117.485 ;
		LAYER VIA3 ;
		RECT 654.555 116.785 654.735 117.485 ;
		LAYER M1 ;
		RECT 654.555 126.045 654.735 126.785 ;
		LAYER M2 ;
		RECT 654.555 126.065 654.735 126.765 ;
		LAYER M3 ;
		RECT 654.555 127.075 654.735 135.035 ;
		LAYER VIA3 ;
		RECT 654.555 127.075 654.735 135.035 ;
		LAYER M3 ;
		RECT 654.555 126.065 654.735 126.765 ;
		LAYER VIA3 ;
		RECT 654.555 126.065 654.735 126.765 ;
		LAYER M3 ;
		RECT 654.555 117.795 654.735 125.755 ;
		LAYER VIA3 ;
		RECT 654.555 117.795 654.735 125.755 ;
		LAYER M2 ;
		RECT 654.555 117.795 654.735 125.755 ;
		LAYER M2 ;
		RECT 654.555 110.835 654.735 116.475 ;
		LAYER M3 ;
		RECT 654.555 110.835 654.735 116.475 ;
		LAYER VIA3 ;
		RECT 654.555 110.835 654.735 116.475 ;
		LAYER M1 ;
		RECT 654.555 172.445 654.735 173.185 ;
		LAYER M2 ;
		RECT 654.555 172.465 654.735 173.165 ;
		LAYER M1 ;
		RECT 654.555 154.895 654.735 162.895 ;
		LAYER M3 ;
		RECT 654.555 172.465 654.735 173.165 ;
		LAYER VIA3 ;
		RECT 654.555 172.465 654.735 173.165 ;
		LAYER M1 ;
		RECT 654.555 164.175 654.735 172.175 ;
		LAYER M3 ;
		RECT 654.555 164.195 654.735 172.155 ;
		LAYER VIA3 ;
		RECT 654.555 164.195 654.735 172.155 ;
		LAYER M2 ;
		RECT 654.555 164.195 654.735 172.155 ;
		LAYER M2 ;
		RECT 654.555 163.185 654.735 163.885 ;
		LAYER M3 ;
		RECT 654.555 163.185 654.735 163.885 ;
		LAYER VIA3 ;
		RECT 654.555 163.185 654.735 163.885 ;
		LAYER M2 ;
		RECT 654.555 153.905 654.735 154.605 ;
		LAYER M3 ;
		RECT 654.555 153.905 654.735 154.605 ;
		LAYER VIA3 ;
		RECT 654.555 153.905 654.735 154.605 ;
		LAYER M1 ;
		RECT 654.555 153.885 654.735 154.625 ;
		LAYER M1 ;
		RECT 654.555 163.165 654.735 163.905 ;
		LAYER M2 ;
		RECT 654.555 154.915 654.735 162.875 ;
		LAYER VIA3 ;
		RECT 654.555 154.915 654.735 162.875 ;
		LAYER M3 ;
		RECT 654.555 154.915 654.735 162.875 ;
		LAYER M1 ;
		RECT 654.555 76.445 654.735 77.185 ;
		LAYER M2 ;
		RECT 654.555 76.465 654.735 77.165 ;
		LAYER M3 ;
		RECT 654.555 76.465 654.735 77.165 ;
		LAYER VIA3 ;
		RECT 654.555 76.465 654.735 77.165 ;
		LAYER M4 ;
		RECT 637.535 80.905 654.735 83.755 ;
		LAYER M4 ;
		RECT 637.535 77.125 654.735 79.115 ;
		LAYER M3 ;
		RECT 654.555 72.835 654.735 76.155 ;
		LAYER VIA3 ;
		RECT 654.555 72.835 654.735 76.155 ;
		LAYER VIA3 ;
		RECT 654.555 63.555 654.735 71.515 ;
		LAYER M1 ;
		RECT 654.555 63.535 654.735 71.535 ;
		LAYER M2 ;
		RECT 654.555 71.825 654.735 72.525 ;
		LAYER M2 ;
		RECT 654.555 17.155 654.735 25.115 ;
		LAYER M3 ;
		RECT 654.555 17.155 654.735 25.115 ;
		LAYER M2 ;
		RECT 654.555 7.875 654.735 15.835 ;
		LAYER M3 ;
		RECT 654.555 7.875 654.735 15.835 ;
		LAYER VIA3 ;
		RECT 654.555 7.875 654.735 15.835 ;
		LAYER M4 ;
		RECT 637.535 59.510 654.345 60.555 ;
		LAYER M4 ;
		RECT 637.535 50.230 654.345 51.275 ;
		LAYER M4 ;
		RECT 637.535 43.785 654.345 44.780 ;
		LAYER M4 ;
		RECT 637.535 40.950 654.345 41.995 ;
		LAYER M4 ;
		RECT 637.535 53.065 654.345 54.060 ;
		LAYER M4 ;
		RECT 637.535 71.625 654.345 72.620 ;
		LAYER M1 ;
		RECT 654.555 72.815 654.735 76.175 ;
		LAYER M2 ;
		RECT 654.555 72.835 654.735 76.155 ;
		LAYER M4 ;
		RECT 637.535 68.790 654.345 69.835 ;
		LAYER M4 ;
		RECT 637.535 62.345 654.345 63.340 ;
		LAYER M4 ;
		RECT 637.535 25.225 654.345 26.220 ;
		LAYER M4 ;
		RECT 637.535 22.390 654.345 23.435 ;
		LAYER M4 ;
		RECT 637.535 15.945 654.345 16.940 ;
		LAYER M4 ;
		RECT 637.535 13.110 654.345 14.155 ;
		LAYER M4 ;
		RECT 637.535 172.265 654.345 173.260 ;
		LAYER M4 ;
		RECT 637.535 169.430 654.345 170.475 ;
		LAYER M4 ;
		RECT 637.535 153.705 654.345 154.700 ;
		LAYER M4 ;
		RECT 637.535 160.150 654.345 161.195 ;
		LAYER M4 ;
		RECT 637.535 162.985 654.345 163.980 ;
		LAYER M4 ;
		RECT 637.535 150.870 654.345 151.915 ;
		LAYER M1 ;
		RECT 654.555 135.325 654.735 136.065 ;
		LAYER M3 ;
		RECT 654.555 136.355 654.735 144.315 ;
		LAYER M2 ;
		RECT 654.555 136.355 654.735 144.315 ;
		LAYER M1 ;
		RECT 654.555 136.335 654.735 144.335 ;
		LAYER M4 ;
		RECT 637.535 102.010 654.345 105.515 ;
		LAYER M4 ;
		RECT 637.535 107.305 654.735 110.155 ;
		LAYER M4 ;
		RECT 637.535 132.310 654.345 133.355 ;
		LAYER M4 ;
		RECT 637.535 113.750 654.345 114.795 ;
		LAYER M4 ;
		RECT 637.535 123.030 654.345 124.075 ;
		LAYER M4 ;
		RECT 637.535 116.585 654.345 117.580 ;
		LAYER M4 ;
		RECT 637.535 141.590 654.345 142.635 ;
		LAYER M4 ;
		RECT 637.535 144.425 654.345 145.420 ;
		LAYER M4 ;
		RECT 637.535 135.145 654.345 136.140 ;
		LAYER M1 ;
		RECT 654.555 173.455 654.735 181.455 ;
		LAYER M2 ;
		RECT 654.555 173.475 654.735 181.435 ;
		LAYER M3 ;
		RECT 654.555 173.475 654.735 181.435 ;
		LAYER VIA3 ;
		RECT 654.555 173.475 654.735 181.435 ;
		LAYER M4 ;
		RECT 637.535 181.545 654.345 182.540 ;
		LAYER VIA3 ;
		RECT 654.555 181.745 654.735 182.445 ;
		LAYER M1 ;
		RECT 654.555 181.725 654.735 182.465 ;
		LAYER M4 ;
		RECT 637.535 178.710 654.345 179.755 ;
		LAYER M4 ;
		RECT 565.275 181.545 637.535 182.040 ;
		LAYER M4 ;
		RECT 565.275 172.265 637.535 172.760 ;
		LAYER M4 ;
		RECT 548.045 176.150 565.275 178.030 ;
		LAYER M4 ;
		RECT 548.045 162.985 565.275 163.515 ;
		LAYER M4 ;
		RECT 548.045 161.055 565.275 161.195 ;
		LAYER M4 ;
		RECT 548.045 157.590 565.275 159.470 ;
		LAYER M4 ;
		RECT 548.045 155.380 565.275 157.425 ;
		LAYER M4 ;
		RECT 565.275 162.985 637.535 163.480 ;
		LAYER M4 ;
		RECT 548.045 56.950 565.275 58.830 ;
		LAYER M4 ;
		RECT 548.045 73.300 565.275 75.345 ;
		LAYER M4 ;
		RECT 548.045 69.695 565.275 69.835 ;
		LAYER M4 ;
		RECT 548.045 60.415 565.275 60.555 ;
		LAYER M4 ;
		RECT 548.045 64.020 565.275 66.065 ;
		LAYER M4 ;
		RECT 548.045 78.975 565.275 79.115 ;
		LAYER M4 ;
		RECT 548.045 80.905 565.275 81.435 ;
		LAYER M4 ;
		RECT 548.045 82.580 565.275 84.625 ;
		LAYER M4 ;
		RECT 548.045 75.510 565.275 77.390 ;
		LAYER M4 ;
		RECT 548.045 54.740 565.275 56.785 ;
		LAYER M4 ;
		RECT 548.045 53.065 565.275 53.595 ;
		LAYER M4 ;
		RECT 548.045 101.910 565.275 103.790 ;
		LAYER M4 ;
		RECT 548.045 111.190 565.275 113.070 ;
		LAYER M4 ;
		RECT 548.045 108.980 565.275 111.025 ;
		LAYER M4 ;
		RECT 548.045 107.305 565.275 107.835 ;
		LAYER M4 ;
		RECT 548.045 105.375 565.275 105.515 ;
		LAYER M4 ;
		RECT 548.045 25.225 565.275 25.755 ;
		LAYER M4 ;
		RECT 548.045 23.295 565.275 23.435 ;
		LAYER M4 ;
		RECT 548.045 10.550 565.275 12.430 ;
		LAYER M4 ;
		RECT 565.275 43.785 637.535 44.280 ;
		LAYER M4 ;
		RECT 548.045 38.390 565.275 40.270 ;
		LAYER M4 ;
		RECT 565.275 25.225 637.535 25.720 ;
		LAYER M4 ;
		RECT 565.275 34.505 637.535 35.000 ;
		LAYER M4 ;
		RECT 565.275 53.065 637.535 53.560 ;
		LAYER M4 ;
		RECT 565.275 71.625 637.535 72.120 ;
		LAYER M4 ;
		RECT 548.045 71.625 565.275 72.155 ;
		LAYER M4 ;
		RECT 565.275 80.905 637.535 81.400 ;
		LAYER M4 ;
		RECT 565.275 107.305 637.535 107.800 ;
		LAYER M4 ;
		RECT 548.045 62.345 565.275 62.875 ;
		LAYER M4 ;
		RECT 548.045 66.230 565.275 68.110 ;
		LAYER M4 ;
		RECT 565.275 125.865 637.535 126.360 ;
		LAYER M4 ;
		RECT 565.275 116.585 637.535 117.080 ;
		LAYER M4 ;
		RECT 565.275 62.345 637.535 62.840 ;
		LAYER M4 ;
		RECT 548.045 26.900 565.275 28.945 ;
		LAYER M4 ;
		RECT 548.045 32.575 565.275 32.715 ;
		LAYER M4 ;
		RECT 548.045 34.505 565.275 35.035 ;
		LAYER M4 ;
		RECT 548.045 36.180 565.275 38.225 ;
		LAYER M4 ;
		RECT 548.045 29.110 565.275 30.990 ;
		LAYER M4 ;
		RECT 548.045 17.620 565.275 19.665 ;
		LAYER M4 ;
		RECT 548.045 15.945 565.275 16.475 ;
		LAYER M4 ;
		RECT 548.045 14.015 565.275 14.155 ;
		LAYER M4 ;
		RECT 548.045 19.830 565.275 21.710 ;
		LAYER M4 ;
		RECT 565.275 6.665 637.535 7.160 ;
		LAYER M4 ;
		RECT 565.275 15.945 637.535 16.440 ;
		LAYER M4 ;
		RECT 548.045 4.735 565.275 4.875 ;
		LAYER M4 ;
		RECT 548.045 1.270 565.275 3.150 ;
		LAYER M4 ;
		RECT 548.045 6.665 565.275 7.195 ;
		LAYER M4 ;
		RECT 548.045 8.340 565.275 10.385 ;
		LAYER M4 ;
		RECT 637.535 6.665 654.345 7.660 ;
		LAYER M4 ;
		RECT 637.535 3.830 654.345 4.875 ;
		LAYER M4 ;
		RECT 637.535 31.670 654.345 32.715 ;
		LAYER M4 ;
		RECT 637.535 34.505 654.345 35.500 ;
		LAYER M1 ;
		RECT 654.555 7.855 654.735 15.855 ;
		LAYER M1 ;
		RECT 654.555 6.845 654.735 7.585 ;
		LAYER M4 ;
		RECT 637.535 125.865 654.345 126.860 ;
		LAYER M4 ;
		RECT 635.910 93.025 654.735 93.385 ;
		LAYER M4 ;
		RECT 548.045 136.820 565.275 138.865 ;
		LAYER M4 ;
		RECT 548.045 135.145 565.275 135.675 ;
		LAYER M4 ;
		RECT 565.275 135.145 637.535 135.640 ;
		LAYER M4 ;
		RECT 548.045 51.135 565.275 51.275 ;
		LAYER M4 ;
		RECT 548.045 47.670 565.275 49.550 ;
		LAYER M4 ;
		RECT 548.045 41.855 565.275 41.995 ;
		LAYER M4 ;
		RECT 548.045 45.460 565.275 47.505 ;
		LAYER M4 ;
		RECT 548.045 43.785 565.275 44.315 ;
		LAYER M4 ;
		RECT 548.045 133.215 565.275 133.355 ;
		LAYER M4 ;
		RECT 548.045 139.030 565.275 140.910 ;
		LAYER M4 ;
		RECT 548.045 142.495 565.275 142.635 ;
		LAYER M4 ;
		RECT 548.045 129.750 565.275 131.630 ;
		LAYER M4 ;
		RECT 548.045 127.540 565.275 129.585 ;
		LAYER M4 ;
		RECT 548.045 125.865 565.275 126.395 ;
		LAYER M4 ;
		RECT 548.045 123.935 565.275 124.075 ;
		LAYER M4 ;
		RECT 548.045 114.655 565.275 114.795 ;
		LAYER M4 ;
		RECT 548.045 116.585 565.275 117.115 ;
		LAYER M4 ;
		RECT 548.045 118.260 565.275 120.305 ;
		LAYER M4 ;
		RECT 548.045 120.470 565.275 122.350 ;
		LAYER M4 ;
		RECT 548.045 179.615 565.275 179.755 ;
		LAYER M4 ;
		RECT 548.045 172.265 565.275 172.795 ;
		LAYER M4 ;
		RECT 548.045 170.335 565.275 170.475 ;
		LAYER M4 ;
		RECT 548.045 166.870 565.275 168.750 ;
		LAYER M4 ;
		RECT 548.045 164.660 565.275 166.705 ;
		LAYER M4 ;
		RECT 548.045 173.940 565.275 175.985 ;
		LAYER M4 ;
		RECT 548.045 153.705 565.275 154.235 ;
		LAYER M4 ;
		RECT 548.045 151.775 565.275 151.915 ;
		LAYER M4 ;
		RECT 548.045 148.310 565.275 150.190 ;
		LAYER M4 ;
		RECT 548.045 146.100 565.275 148.145 ;
		LAYER M4 ;
		RECT 565.275 153.705 637.535 154.200 ;
		LAYER M4 ;
		RECT 548.045 144.425 565.275 144.955 ;
		LAYER M4 ;
		RECT 565.275 144.425 637.535 144.920 ;
		LAYER M4 ;
		RECT 71.735 170.335 88.965 170.475 ;
		LAYER M4 ;
		RECT 71.735 6.665 88.965 7.195 ;
		LAYER M4 ;
		RECT 71.735 1.270 88.965 3.150 ;
		LAYER M4 ;
		RECT 71.735 4.735 88.965 4.875 ;
		LAYER M4 ;
		RECT 71.735 142.495 88.965 142.635 ;
		LAYER M4 ;
		RECT 71.735 139.030 88.965 140.910 ;
		LAYER M4 ;
		RECT 71.735 135.145 88.965 135.675 ;
		LAYER M4 ;
		RECT 71.735 127.540 88.965 129.585 ;
		LAYER M4 ;
		RECT 71.735 133.215 88.965 133.355 ;
		LAYER M4 ;
		RECT 71.735 82.580 88.965 84.625 ;
		LAYER M4 ;
		RECT 71.735 78.975 88.965 79.115 ;
		LAYER M4 ;
		RECT 71.735 75.510 88.965 77.390 ;
		LAYER M4 ;
		RECT 71.735 62.345 88.965 62.875 ;
		LAYER M4 ;
		RECT 71.735 64.020 88.965 66.065 ;
		LAYER M4 ;
		RECT 71.735 80.905 88.965 81.435 ;
		LAYER M4 ;
		RECT 71.735 144.425 88.965 144.955 ;
		LAYER M4 ;
		RECT 71.735 120.470 88.965 122.350 ;
		LAYER M4 ;
		RECT 71.735 125.865 88.965 126.395 ;
		LAYER M4 ;
		RECT 71.735 164.660 88.965 166.705 ;
		LAYER M4 ;
		RECT 71.735 162.985 88.965 163.515 ;
		LAYER M4 ;
		RECT 71.735 151.775 88.965 151.915 ;
		LAYER M4 ;
		RECT 71.735 166.870 88.965 168.750 ;
		LAYER M4 ;
		RECT 71.735 108.980 88.965 111.025 ;
		LAYER M4 ;
		RECT 71.735 101.910 88.965 103.790 ;
		LAYER M4 ;
		RECT 71.735 123.935 88.965 124.075 ;
		LAYER M4 ;
		RECT 71.735 129.750 88.965 131.630 ;
		LAYER M4 ;
		RECT 71.735 105.375 88.965 105.515 ;
		LAYER M4 ;
		RECT 71.735 148.310 88.965 150.190 ;
		LAYER M4 ;
		RECT 71.735 146.100 88.965 148.145 ;
		LAYER M4 ;
		RECT 71.735 136.820 88.965 138.865 ;
		LAYER M4 ;
		RECT 71.735 118.260 88.965 120.305 ;
		LAYER M4 ;
		RECT 71.735 116.585 88.965 117.115 ;
		LAYER M4 ;
		RECT 71.735 114.655 88.965 114.795 ;
		LAYER M4 ;
		RECT 71.735 111.190 88.965 113.070 ;
		LAYER M4 ;
		RECT 71.735 157.590 88.965 159.470 ;
		LAYER M4 ;
		RECT 71.735 161.055 88.965 161.195 ;
		LAYER M4 ;
		RECT 71.735 155.380 88.965 157.425 ;
		LAYER M4 ;
		RECT 71.735 153.705 88.965 154.235 ;
		LAYER M4 ;
		RECT 230.505 155.380 247.735 157.425 ;
		LAYER M4 ;
		RECT 230.505 133.215 247.735 133.355 ;
		LAYER M4 ;
		RECT 230.505 151.775 247.735 151.915 ;
		LAYER M4 ;
		RECT 230.505 127.540 247.735 129.585 ;
		LAYER M4 ;
		RECT 230.505 125.865 247.735 126.395 ;
		LAYER M4 ;
		RECT 230.505 142.495 247.735 142.635 ;
		LAYER M4 ;
		RECT 230.505 139.030 247.735 140.910 ;
		LAYER M4 ;
		RECT 230.505 136.820 247.735 138.865 ;
		LAYER M4 ;
		RECT 230.505 135.145 247.735 135.675 ;
		LAYER M4 ;
		RECT 230.505 64.020 247.735 66.065 ;
		LAYER M4 ;
		RECT 88.965 71.625 230.505 72.120 ;
		LAYER M4 ;
		RECT 88.965 53.065 230.505 53.560 ;
		LAYER M4 ;
		RECT 88.965 43.785 230.505 44.280 ;
		LAYER M4 ;
		RECT 88.965 62.345 230.505 62.840 ;
		LAYER M4 ;
		RECT 160.085 100.005 229.905 100.585 ;
		LAYER M4 ;
		RECT 88.965 125.865 230.505 126.360 ;
		LAYER M4 ;
		RECT 88.965 116.585 230.505 117.080 ;
		LAYER M4 ;
		RECT 160.085 100.585 194.645 101.540 ;
		LAYER M4 ;
		RECT 88.965 107.305 230.505 107.800 ;
		LAYER M4 ;
		RECT 195.345 100.585 229.905 101.540 ;
		LAYER M4 ;
		RECT 88.965 15.945 230.505 16.440 ;
		LAYER M4 ;
		RECT 88.965 6.665 230.505 7.160 ;
		LAYER M4 ;
		RECT 88.965 34.505 230.505 35.000 ;
		LAYER M4 ;
		RECT 88.965 25.225 230.505 25.720 ;
		LAYER M4 ;
		RECT 88.965 144.425 230.505 144.920 ;
		LAYER M4 ;
		RECT 88.965 162.985 230.505 163.480 ;
		LAYER M4 ;
		RECT 88.965 135.145 230.505 135.640 ;
		LAYER M4 ;
		RECT 88.965 153.705 230.505 154.200 ;
		LAYER M4 ;
		RECT 230.505 114.655 247.735 114.795 ;
		LAYER M4 ;
		RECT 230.505 116.585 247.735 117.115 ;
		LAYER M4 ;
		RECT 230.505 118.260 247.735 120.305 ;
		LAYER M4 ;
		RECT 230.505 129.750 247.735 131.630 ;
		LAYER M4 ;
		RECT 230.505 108.980 247.735 111.025 ;
		LAYER M4 ;
		RECT 230.505 107.305 247.735 107.835 ;
		LAYER M4 ;
		RECT 230.505 105.375 247.735 105.515 ;
		LAYER M4 ;
		RECT 230.505 111.190 247.735 113.070 ;
		LAYER M4 ;
		RECT 230.505 10.550 247.735 12.430 ;
		LAYER M4 ;
		RECT 230.505 4.735 247.735 4.875 ;
		LAYER M4 ;
		RECT 230.505 1.270 247.735 3.150 ;
		LAYER M4 ;
		RECT 230.505 8.340 247.735 10.385 ;
		LAYER M4 ;
		RECT 230.505 6.665 247.735 7.195 ;
		LAYER M4 ;
		RECT 230.505 170.335 247.735 170.475 ;
		LAYER M4 ;
		RECT 230.505 146.100 247.735 148.145 ;
		LAYER M4 ;
		RECT 230.505 148.310 247.735 150.190 ;
		LAYER M4 ;
		RECT 230.505 144.425 247.735 144.955 ;
		LAYER M4 ;
		RECT 230.505 157.590 247.735 159.470 ;
		LAYER M4 ;
		RECT 230.505 153.705 247.735 154.235 ;
		LAYER M4 ;
		RECT 230.505 82.580 247.735 84.625 ;
		LAYER M4 ;
		RECT 230.505 80.905 247.735 81.435 ;
		LAYER M4 ;
		RECT 230.505 78.975 247.735 79.115 ;
		LAYER M4 ;
		RECT 230.505 69.695 247.735 69.835 ;
		LAYER M4 ;
		RECT 230.505 73.300 247.735 75.345 ;
		LAYER M4 ;
		RECT 230.505 71.625 247.735 72.155 ;
		LAYER M4 ;
		RECT 230.505 101.910 247.735 103.790 ;
		LAYER M4 ;
		RECT 230.505 54.740 247.735 56.785 ;
		LAYER M4 ;
		RECT 230.505 53.065 247.735 53.595 ;
		LAYER M4 ;
		RECT 230.505 45.460 247.735 47.505 ;
		LAYER M4 ;
		RECT 230.505 25.225 247.735 25.755 ;
		LAYER M4 ;
		RECT 230.505 23.295 247.735 23.435 ;
		LAYER M4 ;
		RECT 230.505 29.110 247.735 30.990 ;
		LAYER M4 ;
		RECT 230.505 26.900 247.735 28.945 ;
		LAYER M4 ;
		RECT 230.505 47.670 247.735 49.550 ;
		LAYER M4 ;
		RECT 230.505 14.015 247.735 14.155 ;
		LAYER M4 ;
		RECT 230.505 17.620 247.735 19.665 ;
		LAYER M4 ;
		RECT 230.505 15.945 247.735 16.475 ;
		LAYER M4 ;
		RECT 230.505 51.135 247.735 51.275 ;
		LAYER M4 ;
		RECT 230.505 19.830 247.735 21.710 ;
		LAYER M4 ;
		RECT 230.505 43.785 247.735 44.315 ;
		LAYER M4 ;
		RECT 230.505 38.390 247.735 40.270 ;
		LAYER M4 ;
		RECT 230.505 36.180 247.735 38.225 ;
		LAYER M4 ;
		RECT 230.505 32.575 247.735 32.715 ;
		LAYER M4 ;
		RECT 230.505 34.505 247.735 35.035 ;
		LAYER M4 ;
		RECT 230.505 66.230 247.735 68.110 ;
		LAYER M4 ;
		RECT 230.505 62.345 247.735 62.875 ;
		LAYER M4 ;
		RECT 230.505 60.415 247.735 60.555 ;
		LAYER M4 ;
		RECT 230.505 56.950 247.735 58.830 ;
		LAYER M4 ;
		RECT 71.735 53.065 88.965 53.595 ;
		LAYER M4 ;
		RECT 71.735 66.230 88.965 68.110 ;
		LAYER M4 ;
		RECT 71.735 71.625 88.965 72.155 ;
		LAYER M4 ;
		RECT 71.735 73.300 88.965 75.345 ;
		LAYER M4 ;
		RECT 71.735 69.695 88.965 69.835 ;
		LAYER M4 ;
		RECT 71.735 26.900 88.965 28.945 ;
		LAYER M4 ;
		RECT 71.735 19.830 88.965 21.710 ;
		LAYER M4 ;
		RECT 71.735 17.620 88.965 19.665 ;
		LAYER M4 ;
		RECT 71.735 15.945 88.965 16.475 ;
		LAYER M4 ;
		RECT 71.735 23.295 88.965 23.435 ;
		LAYER M4 ;
		RECT 71.735 25.225 88.965 25.755 ;
		LAYER M4 ;
		RECT 71.735 38.390 88.965 40.270 ;
		LAYER M4 ;
		RECT 71.735 36.180 88.965 38.225 ;
		LAYER M4 ;
		RECT 71.735 34.505 88.965 35.035 ;
		LAYER M4 ;
		RECT 71.735 32.575 88.965 32.715 ;
		LAYER M4 ;
		RECT 71.735 43.785 88.965 44.315 ;
		LAYER M4 ;
		RECT 71.735 8.340 88.965 10.385 ;
		LAYER M4 ;
		RECT 71.735 10.550 88.965 12.430 ;
		LAYER M4 ;
		RECT 71.735 51.135 88.965 51.275 ;
		LAYER M4 ;
		RECT 71.735 47.670 88.965 49.550 ;
		LAYER M4 ;
		RECT 71.735 45.460 88.965 47.505 ;
		LAYER M4 ;
		RECT 71.735 41.855 88.965 41.995 ;
		LAYER M4 ;
		RECT 71.735 14.015 88.965 14.155 ;
		LAYER M4 ;
		RECT 71.735 29.110 88.965 30.990 ;
		LAYER M4 ;
		RECT 389.275 123.935 406.505 124.075 ;
		LAYER M4 ;
		RECT 389.275 120.470 406.505 122.350 ;
		LAYER M4 ;
		RECT 389.275 116.585 406.505 117.115 ;
		LAYER M4 ;
		RECT 389.275 114.655 406.505 114.795 ;
		LAYER M4 ;
		RECT 389.275 125.865 406.505 126.395 ;
		LAYER M4 ;
		RECT 389.275 133.215 406.505 133.355 ;
		LAYER M4 ;
		RECT 389.275 111.190 406.505 113.070 ;
		LAYER M4 ;
		RECT 389.275 54.740 406.505 56.785 ;
		LAYER M4 ;
		RECT 389.275 56.950 406.505 58.830 ;
		LAYER M4 ;
		RECT 389.275 78.975 406.505 79.115 ;
		LAYER M4 ;
		RECT 389.275 82.580 406.505 84.625 ;
		LAYER M4 ;
		RECT 0.000 172.265 71.735 172.760 ;
		LAYER M4 ;
		RECT 71.735 173.940 88.965 175.985 ;
		LAYER M4 ;
		RECT 71.735 176.150 88.965 178.030 ;
		LAYER M4 ;
		RECT 0.000 179.615 1.365 179.755 ;
		LAYER M4 ;
		RECT 71.735 179.615 88.965 179.755 ;
		LAYER M4 ;
		RECT 71.735 172.265 88.965 172.795 ;
		LAYER M4 ;
		RECT 230.505 164.660 247.735 166.705 ;
		LAYER M4 ;
		RECT 230.505 166.870 247.735 168.750 ;
		LAYER M4 ;
		RECT 230.505 173.940 247.735 175.985 ;
		LAYER M4 ;
		RECT 230.505 176.150 247.735 178.030 ;
		LAYER M4 ;
		RECT 230.505 162.985 247.735 163.515 ;
		LAYER M4 ;
		RECT 230.505 161.055 247.735 161.195 ;
		LAYER M4 ;
		RECT 230.505 179.615 247.735 179.755 ;
		LAYER M4 ;
		RECT 247.735 172.265 389.275 172.760 ;
		LAYER M4 ;
		RECT 230.505 172.265 247.735 172.795 ;
		LAYER M4 ;
		RECT 0.000 170.805 654.345 171.885 ;
		LAYER M4 ;
		RECT 247.735 162.985 389.275 163.480 ;
		LAYER M4 ;
		RECT 0.000 162.985 71.735 163.480 ;
		LAYER M4 ;
		RECT 88.965 172.265 230.505 172.760 ;
		LAYER M4 ;
		RECT 548.045 181.545 565.275 182.075 ;
		LAYER M4 ;
		RECT 406.505 181.545 548.045 182.040 ;
		LAYER M4 ;
		RECT 389.275 181.545 406.505 182.075 ;
		LAYER M4 ;
		RECT 247.735 181.545 389.275 182.040 ;
		LAYER M4 ;
		RECT 0.000 180.085 654.345 181.165 ;
		LAYER M4 ;
		RECT 0.000 181.545 71.735 182.040 ;
		LAYER M4 ;
		RECT 230.505 181.545 247.735 182.075 ;
		LAYER M4 ;
		RECT 88.965 181.545 230.505 182.040 ;
		LAYER M4 ;
		RECT 71.735 181.545 88.965 182.075 ;
		LAYER M4 ;
		RECT 406.505 162.985 548.045 163.480 ;
		LAYER M4 ;
		RECT 389.275 164.660 406.505 166.705 ;
		LAYER M4 ;
		RECT 389.275 161.055 406.505 161.195 ;
		LAYER M4 ;
		RECT 389.275 162.985 406.505 163.515 ;
		LAYER M4 ;
		RECT 0.000 161.525 654.345 162.605 ;
		LAYER M4 ;
		RECT 0.000 161.055 1.365 161.195 ;
		LAYER M4 ;
		RECT 318.855 100.585 353.415 101.540 ;
		LAYER M4 ;
		RECT 248.875 100.585 282.895 101.540 ;
		LAYER M4 ;
		RECT 229.905 100.005 248.335 101.540 ;
		LAYER M4 ;
		RECT 159.385 100.005 160.085 101.540 ;
		LAYER M4 ;
		RECT 36.575 100.585 71.135 101.540 ;
		LAYER M4 ;
		RECT 90.105 100.585 124.125 101.540 ;
		LAYER M4 ;
		RECT 124.825 100.585 159.385 101.540 ;
		LAYER M4 ;
		RECT 89.565 100.005 159.385 100.585 ;
		LAYER M4 ;
		RECT 247.735 135.145 389.275 135.640 ;
		LAYER M4 ;
		RECT 247.735 144.425 389.275 144.920 ;
		LAYER M4 ;
		RECT 230.505 183.220 247.735 185.265 ;
		LAYER M4 ;
		RECT 71.735 183.220 88.965 185.265 ;
		LAYER M4 ;
		RECT 247.735 153.705 389.275 154.200 ;
		LAYER M4 ;
		RECT 0.000 153.705 71.735 154.200 ;
		LAYER M4 ;
		RECT 0.000 152.245 654.345 153.325 ;
		LAYER M4 ;
		RECT 0.000 151.775 1.365 151.915 ;
		LAYER M4 ;
		RECT 0.000 144.425 71.735 144.920 ;
		LAYER M4 ;
		RECT 0.000 142.965 654.345 144.045 ;
		LAYER M4 ;
		RECT 0.000 133.685 654.345 134.765 ;
		LAYER M4 ;
		RECT 0.000 60.415 1.365 60.555 ;
		LAYER M4 ;
		RECT 0.000 105.375 1.365 105.515 ;
		LAYER M4 ;
		RECT 0.000 125.865 71.735 126.360 ;
		LAYER M4 ;
		RECT 0.000 123.935 1.365 124.075 ;
		LAYER M4 ;
		RECT 1.315 100.005 71.135 100.585 ;
		LAYER M4 ;
		RECT 0.000 51.135 1.365 51.275 ;
		LAYER M4 ;
		RECT 0.000 69.695 1.365 69.835 ;
		LAYER M4 ;
		RECT 0.000 116.585 71.735 117.080 ;
		LAYER M4 ;
		RECT 354.115 100.585 374.095 101.540 ;
		LAYER M4 ;
		RECT 318.855 100.005 374.095 100.585 ;
		LAYER M4 ;
		RECT 247.735 62.345 389.275 62.840 ;
		LAYER M4 ;
		RECT 0.000 60.885 654.345 61.965 ;
		LAYER M4 ;
		RECT 0.000 70.165 654.345 71.245 ;
		LAYER M4 ;
		RECT 0.000 71.625 71.735 72.120 ;
		LAYER M4 ;
		RECT 0.000 80.905 71.735 81.400 ;
		LAYER M4 ;
		RECT 0.000 62.345 71.735 62.840 ;
		LAYER M4 ;
		RECT 0.000 53.065 71.735 53.560 ;
		LAYER M4 ;
		RECT 0.000 107.305 71.735 107.800 ;
		LAYER M4 ;
		RECT 0.000 115.125 654.345 116.205 ;
		LAYER M4 ;
		RECT 0.000 51.605 654.345 52.685 ;
		LAYER M4 ;
		RECT 389.275 60.415 406.505 60.555 ;
		LAYER M4 ;
		RECT 389.275 51.135 406.505 51.275 ;
		LAYER M4 ;
		RECT 389.275 47.670 406.505 49.550 ;
		LAYER M4 ;
		RECT 389.275 41.855 406.505 41.995 ;
		LAYER M4 ;
		RECT 389.275 45.460 406.505 47.505 ;
		LAYER M4 ;
		RECT 389.275 43.785 406.505 44.315 ;
		LAYER M4 ;
		RECT 389.275 34.505 406.505 35.035 ;
		LAYER M4 ;
		RECT 389.275 32.575 406.505 32.715 ;
		LAYER M4 ;
		RECT 389.275 36.180 406.505 38.225 ;
		LAYER M4 ;
		RECT 389.275 38.390 406.505 40.270 ;
		LAYER M4 ;
		RECT 389.275 8.340 406.505 10.385 ;
		LAYER M4 ;
		RECT 389.275 10.550 406.505 12.430 ;
		LAYER M4 ;
		RECT 389.275 15.945 406.505 16.475 ;
		LAYER M4 ;
		RECT 389.275 17.620 406.505 19.665 ;
		LAYER M4 ;
		RECT 389.275 14.015 406.505 14.155 ;
		LAYER M4 ;
		RECT 406.505 53.065 548.045 53.560 ;
		LAYER M4 ;
		RECT 389.275 53.065 406.505 53.595 ;
		LAYER M4 ;
		RECT 406.505 15.945 548.045 16.440 ;
		LAYER M4 ;
		RECT 406.505 43.785 548.045 44.280 ;
		LAYER M4 ;
		RECT 406.505 25.225 548.045 25.720 ;
		LAYER M4 ;
		RECT 406.505 34.505 548.045 35.000 ;
		LAYER M4 ;
		RECT 389.275 6.665 406.505 7.195 ;
		LAYER M4 ;
		RECT 389.275 4.735 406.505 4.875 ;
		LAYER M4 ;
		RECT 389.275 1.270 406.505 3.150 ;
		LAYER M4 ;
		RECT 389.275 26.900 406.505 28.945 ;
		LAYER M4 ;
		RECT 389.275 29.110 406.505 30.990 ;
		LAYER M4 ;
		RECT 389.275 19.830 406.505 21.710 ;
		LAYER M4 ;
		RECT 389.275 25.225 406.505 25.755 ;
		LAYER M4 ;
		RECT 389.275 23.295 406.505 23.435 ;
		LAYER M1 ;
		RECT 654.555 182.735 654.735 186.370 ;
		LAYER M2 ;
		RECT 654.555 182.755 654.735 186.370 ;
		LAYER M3 ;
		RECT 654.555 182.755 654.735 186.370 ;
		LAYER M2 ;
		RECT 654.555 181.745 654.735 182.445 ;
		LAYER VIA3 ;
		RECT 654.555 182.755 654.735 186.370 ;
		LAYER M3 ;
		RECT 654.555 181.745 654.735 182.445 ;
		LAYER M4 ;
		RECT 548.045 183.220 565.275 185.265 ;
		LAYER M4 ;
		RECT 389.275 155.380 406.505 157.425 ;
		LAYER M4 ;
		RECT 406.505 172.265 548.045 172.760 ;
		LAYER M4 ;
		RECT 406.505 144.425 548.045 144.920 ;
		LAYER M4 ;
		RECT 406.505 125.865 548.045 126.360 ;
		LAYER M4 ;
		RECT 406.505 6.665 548.045 7.160 ;
		LAYER M4 ;
		RECT 389.275 183.220 406.505 185.265 ;
		LAYER M4 ;
		RECT 389.275 166.870 406.505 168.750 ;
		LAYER M4 ;
		RECT 389.275 157.590 406.505 159.470 ;
		LAYER M4 ;
		RECT 389.275 179.615 406.505 179.755 ;
		LAYER M4 ;
		RECT 389.275 176.150 406.505 178.030 ;
		LAYER M4 ;
		RECT 389.275 172.265 406.505 172.795 ;
		LAYER M4 ;
		RECT 389.275 170.335 406.505 170.475 ;
		LAYER M4 ;
		RECT 389.275 173.940 406.505 175.985 ;
		LAYER M4 ;
		RECT 406.505 107.305 548.045 107.800 ;
		LAYER M4 ;
		RECT 406.505 80.905 548.045 81.400 ;
		LAYER M4 ;
		RECT 406.505 71.625 548.045 72.120 ;
		LAYER M4 ;
		RECT 406.505 62.345 548.045 62.840 ;
		LAYER M4 ;
		RECT 389.275 151.775 406.505 151.915 ;
		LAYER M4 ;
		RECT 389.275 153.705 406.505 154.235 ;
		LAYER M4 ;
		RECT 389.275 64.020 406.505 66.065 ;
		LAYER M4 ;
		RECT 389.275 62.345 406.505 62.875 ;
		LAYER M4 ;
		RECT 406.505 153.705 548.045 154.200 ;
		LAYER M4 ;
		RECT 389.275 127.540 406.505 129.585 ;
		LAYER M4 ;
		RECT 389.275 118.260 406.505 120.305 ;
		LAYER M4 ;
		RECT 406.505 135.145 548.045 135.640 ;
		LAYER M4 ;
		RECT 406.505 116.585 548.045 117.080 ;
		LAYER M4 ;
		RECT 389.275 148.310 406.505 150.190 ;
		LAYER M4 ;
		RECT 389.275 146.100 406.505 148.145 ;
		LAYER M4 ;
		RECT 389.275 108.980 406.505 111.025 ;
		LAYER M4 ;
		RECT 389.275 144.425 406.505 144.955 ;
		LAYER M4 ;
		RECT 389.275 142.495 406.505 142.635 ;
		LAYER M4 ;
		RECT 389.275 139.030 406.505 140.910 ;
		LAYER M4 ;
		RECT 389.275 129.750 406.505 131.630 ;
		LAYER M4 ;
		RECT 389.275 135.145 406.505 135.675 ;
		LAYER M4 ;
		RECT 389.275 136.820 406.505 138.865 ;
		LAYER M4 ;
		RECT 389.275 80.905 406.505 81.435 ;
		LAYER M4 ;
		RECT 389.275 75.510 406.505 77.390 ;
		LAYER M4 ;
		RECT 389.275 71.625 406.505 72.155 ;
		LAYER M4 ;
		RECT 389.275 69.695 406.505 69.835 ;
		LAYER M4 ;
		RECT 389.275 73.300 406.505 75.345 ;
		LAYER M4 ;
		RECT 389.275 66.230 406.505 68.110 ;
		LAYER M4 ;
		RECT 389.275 101.910 406.505 103.790 ;
		LAYER M4 ;
		RECT 389.275 105.375 406.505 105.515 ;
		LAYER M4 ;
		RECT 389.275 107.305 406.505 107.835 ;
		LAYER M4 ;
		RECT 318.155 100.005 318.855 101.540 ;
		LAYER M4 ;
		RECT 248.335 100.005 318.155 100.585 ;
		LAYER M4 ;
		RECT 247.735 107.305 389.275 107.800 ;
		LAYER M4 ;
		RECT 283.595 100.585 318.155 101.540 ;
		LAYER M4 ;
		RECT 230.505 123.935 247.735 124.075 ;
		LAYER M4 ;
		RECT 230.505 120.470 247.735 122.350 ;
		LAYER M4 ;
		RECT 247.735 125.865 389.275 126.360 ;
		LAYER M4 ;
		RECT 247.735 116.585 389.275 117.080 ;
		LAYER M4 ;
		RECT 247.735 80.905 389.275 81.400 ;
		LAYER M4 ;
		RECT 247.735 71.625 389.275 72.120 ;
		LAYER M4 ;
		RECT 247.735 53.065 389.275 53.560 ;
		LAYER M4 ;
		RECT 247.735 25.225 389.275 25.720 ;
		LAYER M4 ;
		RECT 247.735 43.785 389.275 44.280 ;
		LAYER M4 ;
		RECT 247.735 34.505 389.275 35.000 ;
		LAYER M4 ;
		RECT 230.505 75.510 247.735 77.390 ;
		LAYER M4 ;
		RECT 230.505 41.855 247.735 41.995 ;
		LAYER M4 ;
		RECT 247.735 15.945 389.275 16.440 ;
		LAYER M4 ;
		RECT 71.735 107.305 88.965 107.835 ;
		LAYER M4 ;
		RECT 71.735 60.415 88.965 60.555 ;
		LAYER M4 ;
		RECT 71.735 56.950 88.965 58.830 ;
		LAYER M4 ;
		RECT 71.735 54.740 88.965 56.785 ;
		LAYER M4 ;
		RECT 88.965 80.905 230.505 81.400 ;
		LAYER M4 ;
		RECT 0.000 135.145 71.735 135.640 ;
		LAYER M4 ;
		RECT 0.000 42.325 654.345 43.405 ;
		LAYER M4 ;
		RECT 0.000 43.785 71.735 44.280 ;
		LAYER M4 ;
		RECT 247.735 6.665 389.275 7.160 ;
		LAYER M2 ;
		RECT 0.000 0.000 654.555 186.370 ;
		LAYER M1 ;
		RECT 0.000 0.000 654.555 186.370 ;
		LAYER M4 ;
		RECT 0.000 4.735 1.365 4.875 ;
		LAYER M4 ;
		RECT 0.000 15.945 71.735 16.440 ;
		LAYER M4 ;
		RECT 0.000 25.225 71.735 25.720 ;
		LAYER M4 ;
		RECT 0.000 34.505 71.735 35.000 ;
		LAYER M4 ;
		RECT 0.000 14.015 1.365 14.155 ;
		LAYER M4 ;
		RECT 0.000 6.665 71.735 7.160 ;
		LAYER M4 ;
		RECT 0.000 14.485 654.345 15.565 ;
		LAYER M4 ;
		RECT 0.000 23.765 654.345 24.845 ;
		LAYER M4 ;
		RECT 0.000 33.045 654.345 34.125 ;
		LAYER M3 ;
		RECT 0.000 0.000 654.555 186.370 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 654.555 186.370 ;
		LAYER M4 ;
		RECT 0.000 5.205 654.345 6.285 ;
		LAYER M4 ;
		RECT 0.000 41.855 1.365 41.995 ;
		LAYER M4 ;
		RECT 0.000 32.575 1.365 32.715 ;
		LAYER M4 ;
		RECT 0.000 23.295 1.365 23.435 ;
		LAYER M4 ;
		RECT 0.000 170.335 1.365 170.475 ;
		LAYER M4 ;
		RECT 0.000 114.655 1.365 114.795 ;
		LAYER M4 ;
		RECT 0.000 78.975 1.365 79.115 ;
		LAYER M4 ;
		RECT 0.000 100.005 1.315 101.540 ;
		LAYER M4 ;
		RECT 0.000 142.495 1.365 142.635 ;
		LAYER M4 ;
		RECT 0.000 133.215 1.365 133.355 ;
		LAYER M4 ;
		RECT 374.095 100.005 654.735 101.540 ;
		LAYER M4 ;
		RECT 0.000 105.845 654.735 106.925 ;
		LAYER M4 ;
		RECT 0.000 93.955 654.735 99.435 ;
		LAYER M4 ;
		RECT 0.000 79.445 654.735 80.525 ;
		LAYER M4 ;
		RECT 0.000 84.535 654.735 90.355 ;
		LAYER M4 ;
		RECT 0.000 124.405 654.345 125.485 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 654.735 186.370 ;
		LAYER M4 ;
		RECT 1.315 100.585 35.875 101.540 ;
		LAYER M4 ;
		RECT 71.135 100.005 89.565 101.540 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 654.735 186.370 ;
	END
	# End of OBS

END TS1N28HPCPHVTB32768X18M16SSO

END LIBRARY
