# Created by MC2 : Version 2012.02.00.d on 2024/05/10, 14:04:38

#*********************************************************************************************************************/
# Software       : TSMC MEMORY COMPILER tsn28hpcpd127spsram_2012.02.00.d.180a						*/
# Technology     : TSMC 28nm CMOS LOGIC High Performance Compact Mobile Computing Plus 1P10M HKMG CU_ELK 0.9V				*/
#  Memory Type    : TSMC 28nm High Performance Compact Mobile Computing Plus Single Port SRAM with d127 bit cell HVT periphery */
# Library Name   : ts1n28hpcphvtb32768x9m16sso (user specify : TS1N28HPCPHVTB32768X9M16SSO)				*/
# Library Version: 180a												*/
# Generated Time : 2024/05/10, 14:04:29										*/
#*********************************************************************************************************************/
#															*/
# STATEMENT OF USE													*/
#															*/
# This information contains confidential and proprietary information of TSMC.					*/
# No part of this information may be reproduced, transmitted, transcribed,						*/
# stored in a retrieval system, or translated into any human or computer						*/
# language, in any form or by any means, electronic, mechanical, magnetic,						*/
# optical, chemical, manual, or otherwise, without the prior written permission					*/
# of TSMC. This information was prepared for informational purpose and is for					*/
# use by TSMC's customers only. TSMC reserves the right to make changes in the					*/
# information at any time and without notice.									*/
#															*/
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS1N28HPCPHVTB32768X9M16SSO
	CLASS BLOCK ;
	FOREIGN TS1N28HPCPHVTB32768X9M16SSO 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 654.735 BY 102.850 ;
	SYMMETRY X Y ;
	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 58.550 654.735 58.700 ;
			LAYER M2 ;
			RECT 654.555 58.550 654.735 58.700 ;
			LAYER M1 ;
			RECT 654.555 58.550 654.735 58.700 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[0]

	PIN A[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 48.690 654.735 48.840 ;
			LAYER M1 ;
			RECT 654.555 48.690 654.735 48.840 ;
			LAYER M3 ;
			RECT 654.555 48.690 654.735 48.840 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[10]

	PIN A[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 48.300 654.735 48.450 ;
			LAYER M3 ;
			RECT 654.555 48.300 654.735 48.450 ;
			LAYER M1 ;
			RECT 654.555 48.300 654.735 48.450 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[11]

	PIN A[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 60.990 654.735 61.140 ;
			LAYER M3 ;
			RECT 654.555 60.990 654.735 61.140 ;
			LAYER M2 ;
			RECT 654.555 60.990 654.735 61.140 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[12]

	PIN A[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 60.600 654.735 60.750 ;
			LAYER M3 ;
			RECT 654.555 60.600 654.735 60.750 ;
			LAYER M2 ;
			RECT 654.555 60.600 654.735 60.750 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[13]

	PIN A[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 58.940 654.735 59.090 ;
			LAYER M2 ;
			RECT 654.555 58.940 654.735 59.090 ;
			LAYER M3 ;
			RECT 654.555 58.940 654.735 59.090 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[14]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 56.890 654.735 57.040 ;
			LAYER M2 ;
			RECT 654.555 56.890 654.735 57.040 ;
			LAYER M3 ;
			RECT 654.555 56.890 654.735 57.040 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 56.500 654.735 56.650 ;
			LAYER M2 ;
			RECT 654.555 56.500 654.735 56.650 ;
			LAYER M1 ;
			RECT 654.555 56.500 654.735 56.650 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 46.640 654.735 46.790 ;
			LAYER M3 ;
			RECT 654.555 46.640 654.735 46.790 ;
			LAYER M1 ;
			RECT 654.555 46.640 654.735 46.790 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 52.400 654.735 52.550 ;
			LAYER M3 ;
			RECT 654.555 52.400 654.735 52.550 ;
			LAYER M2 ;
			RECT 654.555 52.400 654.735 52.550 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 50.740 654.735 50.890 ;
			LAYER M3 ;
			RECT 654.555 50.740 654.735 50.890 ;
			LAYER M1 ;
			RECT 654.555 50.740 654.735 50.890 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 50.350 654.735 50.500 ;
			LAYER M2 ;
			RECT 654.555 50.350 654.735 50.500 ;
			LAYER M3 ;
			RECT 654.555 50.350 654.735 50.500 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 54.840 654.735 54.990 ;
			LAYER M2 ;
			RECT 654.555 54.840 654.735 54.990 ;
			LAYER M3 ;
			RECT 654.555 54.840 654.735 54.990 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 54.450 654.735 54.600 ;
			LAYER M3 ;
			RECT 654.555 54.450 654.735 54.600 ;
			LAYER M2 ;
			RECT 654.555 54.450 654.735 54.600 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 52.790 654.735 52.940 ;
			LAYER M2 ;
			RECT 654.555 52.790 654.735 52.940 ;
			LAYER M3 ;
			RECT 654.555 52.790 654.735 52.940 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[9]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 62.650 654.735 62.800 ;
			LAYER M2 ;
			RECT 654.555 62.650 654.735 62.800 ;
			LAYER M1 ;
			RECT 654.555 62.650 654.735 62.800 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.115300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.228300 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.515900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.249900 LAYER M2 ;
		ANTENNAMAXAREACAR 10.191100 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.732500 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 11.091100 LAYER M3 ;
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 63.280 654.735 63.430 ;
			LAYER M2 ;
			RECT 654.555 63.280 654.735 63.430 ;
			LAYER M1 ;
			RECT 654.555 63.280 654.735 63.430 ;
		END
		ANTENNAGATEAREA 2.013900 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 3.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 5.372500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.331500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA1 ;
		ANTENNAGATEAREA 2.013900 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 2.694600 LAYER M2 ;
		ANTENNAMAXAREACAR 33.912400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.292500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.097200 LAYER VIA2 ;
		ANTENNAGATEAREA 2.013900 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 2.754400 LAYER M3 ;
		ANTENNAMAXAREACAR 35.107800 LAYER M3 ;
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 6.635 654.735 6.785 ;
			LAYER M3 ;
			RECT 654.555 6.635 654.735 6.785 ;
			LAYER M1 ;
			RECT 654.555 6.635 654.735 6.785 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 15.915 654.735 16.065 ;
			LAYER M3 ;
			RECT 654.555 15.915 654.735 16.065 ;
			LAYER M2 ;
			RECT 654.555 15.915 654.735 16.065 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 25.195 654.735 25.345 ;
			LAYER M3 ;
			RECT 654.555 25.195 654.735 25.345 ;
			LAYER M2 ;
			RECT 654.555 25.195 654.735 25.345 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 34.475 654.735 34.625 ;
			LAYER M3 ;
			RECT 654.555 34.475 654.735 34.625 ;
			LAYER M2 ;
			RECT 654.555 34.475 654.735 34.625 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 39.115 654.735 39.265 ;
			LAYER M2 ;
			RECT 654.555 39.115 654.735 39.265 ;
			LAYER M1 ;
			RECT 654.555 39.115 654.735 39.265 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 72.475 654.735 72.625 ;
			LAYER M3 ;
			RECT 654.555 72.475 654.735 72.625 ;
			LAYER M2 ;
			RECT 654.555 72.475 654.735 72.625 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 79.435 654.735 79.585 ;
			LAYER M2 ;
			RECT 654.555 79.435 654.735 79.585 ;
			LAYER M1 ;
			RECT 654.555 79.435 654.735 79.585 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 88.715 654.735 88.865 ;
			LAYER M1 ;
			RECT 654.555 88.715 654.735 88.865 ;
			LAYER M2 ;
			RECT 654.555 88.715 654.735 88.865 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 97.995 654.735 98.145 ;
			LAYER M2 ;
			RECT 654.555 97.995 654.735 98.145 ;
			LAYER M1 ;
			RECT 654.555 97.995 654.735 98.145 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[8]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 7.645 654.735 7.795 ;
			LAYER M2 ;
			RECT 654.555 7.645 654.735 7.795 ;
			LAYER M3 ;
			RECT 654.555 7.645 654.735 7.795 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 16.925 654.735 17.075 ;
			LAYER M3 ;
			RECT 654.555 16.925 654.735 17.075 ;
			LAYER M2 ;
			RECT 654.555 16.925 654.735 17.075 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 26.205 654.735 26.355 ;
			LAYER M3 ;
			RECT 654.555 26.205 654.735 26.355 ;
			LAYER M2 ;
			RECT 654.555 26.205 654.735 26.355 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 35.485 654.735 35.635 ;
			LAYER M2 ;
			RECT 654.555 35.485 654.735 35.635 ;
			LAYER M1 ;
			RECT 654.555 35.485 654.735 35.635 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 40.125 654.735 40.275 ;
			LAYER M1 ;
			RECT 654.555 40.125 654.735 40.275 ;
			LAYER M3 ;
			RECT 654.555 40.125 654.735 40.275 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 73.485 654.735 73.635 ;
			LAYER M1 ;
			RECT 654.555 73.485 654.735 73.635 ;
			LAYER M3 ;
			RECT 654.555 73.485 654.735 73.635 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 80.445 654.735 80.595 ;
			LAYER M3 ;
			RECT 654.555 80.445 654.735 80.595 ;
			LAYER M1 ;
			RECT 654.555 80.445 654.735 80.595 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 89.725 654.735 89.875 ;
			LAYER M3 ;
			RECT 654.555 89.725 654.735 89.875 ;
			LAYER M2 ;
			RECT 654.555 89.725 654.735 89.875 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 99.005 654.735 99.155 ;
			LAYER M1 ;
			RECT 654.555 99.005 654.735 99.155 ;
			LAYER M3 ;
			RECT 654.555 99.005 654.735 99.155 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[8]

	PIN SD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 44.025 654.735 44.175 ;
			LAYER M2 ;
			RECT 654.555 44.025 654.735 44.175 ;
			LAYER M3 ;
			RECT 654.555 44.025 654.735 44.175 ;
		END
		ANTENNAGATEAREA 0.051000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.839700 LAYER M1 ;
		ANTENNAMAXAREACAR 9.087800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.585600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.051000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.499900 LAYER M2 ;
		ANTENNAMAXAREACAR 48.990700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.878400 LAYER VIA2 ;
		ANTENNAGATEAREA 0.051000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.590600 LAYER M3 ;
		ANTENNAMAXAREACAR 48.990700 LAYER M3 ;
	END SD

	PIN SLP
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 44.740 654.735 44.890 ;
			LAYER M2 ;
			RECT 654.555 44.740 654.735 44.890 ;
			LAYER M3 ;
			RECT 654.555 44.740 654.735 44.890 ;
		END
		ANTENNAGATEAREA 0.027000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.172400 LAYER M1 ;
		ANTENNAMAXAREACAR 8.260000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.433300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.027000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.269000 LAYER M2 ;
		ANTENNAMAXAREACAR 48.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.027000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.564300 LAYER M3 ;
		ANTENNAMAXAREACAR 48.814800 LAYER M3 ;
	END SLP

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.000 4.875 654.345 5.205 ;
			LAYER M4 ;
			RECT 0.000 14.155 654.345 14.485 ;
			LAYER M4 ;
			RECT 0.000 23.435 654.345 23.765 ;
			LAYER M4 ;
			RECT 0.000 32.715 654.345 33.045 ;
			LAYER M4 ;
			RECT 0.000 41.995 654.735 42.325 ;
			LAYER M4 ;
			RECT 0.000 54.635 654.735 55.205 ;
			LAYER M4 ;
			RECT 0.000 55.335 654.735 55.905 ;
			LAYER M4 ;
			RECT 0.000 62.315 654.735 62.885 ;
			LAYER M4 ;
			RECT 0.000 68.395 654.735 68.725 ;
			LAYER M4 ;
			RECT 0.000 77.675 654.345 78.005 ;
			LAYER M4 ;
			RECT 0.000 86.955 654.345 87.285 ;
			LAYER M4 ;
			RECT 0.000 96.235 654.345 96.565 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.000 6.285 654.345 6.665 ;
			LAYER M4 ;
			RECT 0.000 15.565 654.345 15.945 ;
			LAYER M4 ;
			RECT 0.000 24.845 654.345 25.225 ;
			LAYER M4 ;
			RECT 0.000 34.125 654.345 34.505 ;
			LAYER M4 ;
			RECT 0.000 43.405 654.735 43.785 ;
			LAYER M4 ;
			RECT 0.000 53.235 654.735 53.805 ;
			LAYER M4 ;
			RECT 0.000 53.935 654.735 54.505 ;
			LAYER M4 ;
			RECT 0.000 56.265 654.735 56.835 ;
			LAYER M4 ;
			RECT 0.000 69.805 654.735 70.185 ;
			LAYER M4 ;
			RECT 0.000 79.085 654.345 79.465 ;
			LAYER M4 ;
			RECT 0.000 88.365 654.345 88.745 ;
			LAYER M4 ;
			RECT 0.000 97.645 654.345 98.025 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 46.250 654.735 46.400 ;
			LAYER M1 ;
			RECT 654.555 46.250 654.735 46.400 ;
			LAYER M3 ;
			RECT 654.555 46.250 654.735 46.400 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.445400 LAYER M2 ;
		ANTENNAMAXAREACAR 16.888300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 17.788300 LAYER M3 ;
	END WEB

	OBS
		# Promoted blockages
		LAYER M2 ;
		RECT 654.555 62.880 654.735 63.200 ;
		LAYER M3 ;
		RECT 654.555 62.880 654.735 63.200 ;
		LAYER M3 ;
		RECT 654.555 89.955 654.735 97.915 ;
		LAYER VIA3 ;
		RECT 654.555 62.880 654.735 63.200 ;
		LAYER M1 ;
		RECT 654.555 80.655 654.735 88.655 ;
		LAYER M1 ;
		RECT 654.555 79.645 654.735 80.385 ;
		LAYER M3 ;
		RECT 654.555 80.675 654.735 88.635 ;
		LAYER VIA3 ;
		RECT 654.555 80.675 654.735 88.635 ;
		LAYER M3 ;
		RECT 654.555 79.665 654.735 80.365 ;
		LAYER VIA3 ;
		RECT 654.555 79.665 654.735 80.365 ;
		LAYER M2 ;
		RECT 654.555 79.665 654.735 80.365 ;
		LAYER M2 ;
		RECT 654.555 88.945 654.735 89.645 ;
		LAYER M1 ;
		RECT 654.555 89.935 654.735 97.935 ;
		LAYER M2 ;
		RECT 654.555 98.225 654.735 98.925 ;
		LAYER M1 ;
		RECT 654.555 98.205 654.735 98.945 ;
		LAYER VIA3 ;
		RECT 654.555 89.955 654.735 97.915 ;
		LAYER M3 ;
		RECT 654.555 88.945 654.735 89.645 ;
		LAYER M2 ;
		RECT 654.555 80.675 654.735 88.635 ;
		LAYER M3 ;
		RECT 654.555 99.235 654.735 102.850 ;
		LAYER M1 ;
		RECT 654.555 88.925 654.735 89.665 ;
		LAYER VIA3 ;
		RECT 654.555 88.945 654.735 89.645 ;
		LAYER M2 ;
		RECT 654.555 99.235 654.735 102.850 ;
		LAYER VIA3 ;
		RECT 654.555 99.235 654.735 102.850 ;
		LAYER M1 ;
		RECT 654.555 72.685 654.735 73.425 ;
		LAYER M3 ;
		RECT 654.555 63.510 654.735 72.395 ;
		LAYER M2 ;
		RECT 654.555 63.510 654.735 72.395 ;
		LAYER VIA3 ;
		RECT 654.555 63.510 654.735 72.395 ;
		LAYER M4 ;
		RECT 654.345 65.250 654.735 68.395 ;
		LAYER M2 ;
		RECT 654.555 72.705 654.735 73.405 ;
		LAYER M3 ;
		RECT 654.555 72.705 654.735 73.405 ;
		LAYER VIA3 ;
		RECT 654.555 72.705 654.735 73.405 ;
		LAYER M4 ;
		RECT 637.535 79.465 654.345 80.460 ;
		LAYER M4 ;
		RECT 637.535 64.890 654.345 68.395 ;
		LAYER M2 ;
		RECT 654.555 89.955 654.735 97.915 ;
		LAYER M3 ;
		RECT 654.555 98.225 654.735 98.925 ;
		LAYER VIA3 ;
		RECT 654.555 98.225 654.735 98.925 ;
		LAYER M1 ;
		RECT 654.555 99.215 654.735 102.850 ;
		LAYER M4 ;
		RECT 637.535 98.025 654.345 99.020 ;
		LAYER M4 ;
		RECT 637.535 95.190 654.345 96.235 ;
		LAYER M4 ;
		RECT 637.535 88.745 654.345 89.740 ;
		LAYER M2 ;
		RECT 654.555 60.830 654.735 60.910 ;
		LAYER M3 ;
		RECT 654.555 60.830 654.735 60.910 ;
		LAYER M2 ;
		RECT 654.555 61.220 654.735 62.570 ;
		LAYER M3 ;
		RECT 654.555 61.220 654.735 62.570 ;
		LAYER VIA3 ;
		RECT 654.555 60.830 654.735 60.910 ;
		LAYER VIA3 ;
		RECT 654.555 61.220 654.735 62.570 ;
		LAYER M3 ;
		RECT 654.555 53.020 654.735 54.370 ;
		LAYER M1 ;
		RECT 654.555 62.860 654.735 63.220 ;
		LAYER M1 ;
		RECT 654.555 61.200 654.735 62.590 ;
		LAYER M1 ;
		RECT 654.555 59.150 654.735 60.540 ;
		LAYER M1 ;
		RECT 654.555 60.810 654.735 60.930 ;
		LAYER M1 ;
		RECT 654.555 56.710 654.735 56.830 ;
		LAYER M2 ;
		RECT 654.555 57.120 654.735 58.470 ;
		LAYER M2 ;
		RECT 654.555 55.070 654.735 56.420 ;
		LAYER M2 ;
		RECT 654.555 59.170 654.735 60.520 ;
		LAYER M3 ;
		RECT 654.555 55.070 654.735 56.420 ;
		LAYER M4 ;
		RECT 635.910 55.905 654.735 56.265 ;
		LAYER M2 ;
		RECT 654.555 53.020 654.735 54.370 ;
		LAYER M2 ;
		RECT 654.555 50.580 654.735 50.660 ;
		LAYER M3 ;
		RECT 654.555 50.580 654.735 50.660 ;
		LAYER M1 ;
		RECT 654.555 52.610 654.735 52.730 ;
		LAYER M2 ;
		RECT 654.555 52.630 654.735 52.710 ;
		LAYER M3 ;
		RECT 654.555 52.630 654.735 52.710 ;
		LAYER M1 ;
		RECT 654.555 50.950 654.735 52.340 ;
		LAYER M3 ;
		RECT 654.555 26.435 654.735 34.395 ;
		LAYER M2 ;
		RECT 654.555 26.435 654.735 34.395 ;
		LAYER M1 ;
		RECT 654.555 26.415 654.735 34.415 ;
		LAYER M3 ;
		RECT 654.555 34.705 654.735 35.405 ;
		LAYER M4 ;
		RECT 637.535 6.665 654.345 7.660 ;
		LAYER M4 ;
		RECT 637.535 34.505 654.345 35.500 ;
		LAYER M4 ;
		RECT 637.535 40.005 654.735 41.995 ;
		LAYER M4 ;
		RECT 637.535 43.785 654.735 46.635 ;
		LAYER M4 ;
		RECT 637.535 22.390 654.345 23.435 ;
		LAYER M4 ;
		RECT 637.535 15.945 654.345 16.940 ;
		LAYER M4 ;
		RECT 637.535 13.110 654.345 14.155 ;
		LAYER M4 ;
		RECT 637.535 31.670 654.345 32.715 ;
		LAYER M4 ;
		RECT 637.535 25.225 654.345 26.220 ;
		LAYER M1 ;
		RECT 654.555 39.325 654.735 40.065 ;
		LAYER M2 ;
		RECT 654.555 39.345 654.735 40.045 ;
		LAYER M2 ;
		RECT 654.555 35.715 654.735 39.035 ;
		LAYER M4 ;
		RECT 565.275 34.505 637.535 35.000 ;
		LAYER M4 ;
		RECT 548.045 34.505 565.275 35.035 ;
		LAYER M4 ;
		RECT 548.045 17.620 565.275 19.665 ;
		LAYER M4 ;
		RECT 548.045 19.830 565.275 21.710 ;
		LAYER M4 ;
		RECT 548.045 32.575 565.275 32.715 ;
		LAYER M4 ;
		RECT 548.045 36.180 565.275 38.225 ;
		LAYER M4 ;
		RECT 548.045 15.945 565.275 16.475 ;
		LAYER M4 ;
		RECT 548.045 10.550 565.275 12.430 ;
		LAYER M4 ;
		RECT 548.045 8.340 565.275 10.385 ;
		LAYER M4 ;
		RECT 565.275 15.945 637.535 16.440 ;
		LAYER M4 ;
		RECT 565.275 43.785 637.535 44.280 ;
		LAYER M4 ;
		RECT 637.535 3.830 654.345 4.875 ;
		LAYER M4 ;
		RECT 565.275 6.665 637.535 7.160 ;
		LAYER M4 ;
		RECT 565.275 25.225 637.535 25.720 ;
		LAYER M4 ;
		RECT 548.045 38.390 565.275 40.270 ;
		LAYER M4 ;
		RECT 548.045 41.855 565.275 41.995 ;
		LAYER M4 ;
		RECT 548.045 43.785 565.275 44.315 ;
		LAYER M4 ;
		RECT 548.045 26.900 565.275 28.945 ;
		LAYER M4 ;
		RECT 548.045 25.225 565.275 25.755 ;
		LAYER M4 ;
		RECT 548.045 23.295 565.275 23.435 ;
		LAYER M4 ;
		RECT 548.045 29.110 565.275 30.990 ;
		LAYER M4 ;
		RECT 548.045 6.665 565.275 7.195 ;
		LAYER M4 ;
		RECT 548.045 4.735 565.275 4.875 ;
		LAYER M4 ;
		RECT 548.045 14.015 565.275 14.155 ;
		LAYER M4 ;
		RECT 406.505 15.945 548.045 16.440 ;
		LAYER M4 ;
		RECT 548.045 1.270 565.275 3.150 ;
		LAYER M4 ;
		RECT 247.735 6.665 389.275 7.160 ;
		LAYER M4 ;
		RECT 406.505 6.665 548.045 7.160 ;
		LAYER M4 ;
		RECT 247.735 15.945 389.275 16.440 ;
		LAYER M4 ;
		RECT 230.505 8.340 247.735 10.385 ;
		LAYER M4 ;
		RECT 389.275 8.340 406.505 10.385 ;
		LAYER M4 ;
		RECT 0.000 14.485 654.345 15.565 ;
		LAYER M4 ;
		RECT 389.275 1.270 406.505 3.150 ;
		LAYER M4 ;
		RECT 389.275 4.735 406.505 4.875 ;
		LAYER M4 ;
		RECT 230.505 1.270 247.735 3.150 ;
		LAYER M4 ;
		RECT 230.505 6.665 247.735 7.195 ;
		LAYER M4 ;
		RECT 389.275 6.665 406.505 7.195 ;
		LAYER M4 ;
		RECT 0.000 5.205 654.345 6.285 ;
		LAYER M4 ;
		RECT 230.505 4.735 247.735 4.875 ;
		LAYER M4 ;
		RECT 71.735 1.270 88.965 3.150 ;
		LAYER M4 ;
		RECT 88.965 6.665 230.505 7.160 ;
		LAYER M4 ;
		RECT 0.000 4.735 1.365 4.875 ;
		LAYER M4 ;
		RECT 0.000 6.665 71.735 7.160 ;
		LAYER M4 ;
		RECT 71.735 6.665 88.965 7.195 ;
		LAYER M4 ;
		RECT 71.735 8.340 88.965 10.385 ;
		LAYER M4 ;
		RECT 71.735 4.735 88.965 4.875 ;
		LAYER M1 ;
		RECT 654.555 73.695 654.735 79.375 ;
		LAYER M2 ;
		RECT 654.555 73.715 654.735 79.355 ;
		LAYER M3 ;
		RECT 654.555 73.715 654.735 79.355 ;
		LAYER VIA3 ;
		RECT 654.555 73.715 654.735 79.355 ;
		LAYER M1 ;
		RECT 654.555 63.490 654.735 72.415 ;
		LAYER M4 ;
		RECT 637.535 70.185 654.735 73.035 ;
		LAYER M4 ;
		RECT 637.535 76.630 654.345 77.675 ;
		LAYER M4 ;
		RECT 637.535 85.910 654.345 86.955 ;
		LAYER M4 ;
		RECT 565.275 79.465 637.535 79.960 ;
		LAYER M4 ;
		RECT 374.095 62.885 654.735 64.420 ;
		LAYER M4 ;
		RECT 565.275 70.185 637.535 70.680 ;
		LAYER M4 ;
		RECT 406.505 70.185 548.045 70.680 ;
		LAYER M4 ;
		RECT 548.045 64.790 565.275 66.670 ;
		LAYER M4 ;
		RECT 548.045 68.255 565.275 68.395 ;
		LAYER M4 ;
		RECT 406.505 79.465 548.045 79.960 ;
		LAYER M4 ;
		RECT 406.505 88.745 548.045 89.240 ;
		LAYER M4 ;
		RECT 548.045 88.745 565.275 89.275 ;
		LAYER M4 ;
		RECT 565.275 88.745 637.535 89.240 ;
		LAYER M4 ;
		RECT 406.505 98.025 548.045 98.520 ;
		LAYER M4 ;
		RECT 565.275 98.025 637.535 98.520 ;
		LAYER M4 ;
		RECT 389.275 34.505 406.505 35.035 ;
		LAYER M4 ;
		RECT 389.275 29.110 406.505 30.990 ;
		LAYER M4 ;
		RECT 389.275 26.900 406.505 28.945 ;
		LAYER M4 ;
		RECT 389.275 25.225 406.505 25.755 ;
		LAYER M4 ;
		RECT 406.505 25.225 548.045 25.720 ;
		LAYER M4 ;
		RECT 406.505 34.505 548.045 35.000 ;
		LAYER M4 ;
		RECT 389.275 36.180 406.505 38.225 ;
		LAYER M4 ;
		RECT 389.275 23.295 406.505 23.435 ;
		LAYER M4 ;
		RECT 389.275 19.830 406.505 21.710 ;
		LAYER M4 ;
		RECT 389.275 14.015 406.505 14.155 ;
		LAYER M4 ;
		RECT 0.000 23.765 654.345 24.845 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 654.735 102.850 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 654.735 102.850 ;
		LAYER M4 ;
		RECT 548.045 70.185 565.275 70.715 ;
		LAYER M4 ;
		RECT 548.045 99.700 565.275 101.745 ;
		LAYER M4 ;
		RECT 548.045 98.025 565.275 98.555 ;
		LAYER M4 ;
		RECT 548.045 77.535 565.275 77.675 ;
		LAYER M4 ;
		RECT 548.045 74.070 565.275 75.950 ;
		LAYER M4 ;
		RECT 548.045 71.860 565.275 73.905 ;
		LAYER M4 ;
		RECT 548.045 86.815 565.275 86.955 ;
		LAYER M4 ;
		RECT 548.045 90.420 565.275 92.465 ;
		LAYER M4 ;
		RECT 548.045 92.630 565.275 94.510 ;
		LAYER M4 ;
		RECT 548.045 96.095 565.275 96.235 ;
		LAYER M4 ;
		RECT 548.045 83.350 565.275 85.230 ;
		LAYER M4 ;
		RECT 548.045 81.140 565.275 83.185 ;
		LAYER M4 ;
		RECT 548.045 79.465 565.275 79.995 ;
		LAYER M4 ;
		RECT 71.735 41.855 88.965 41.995 ;
		LAYER M4 ;
		RECT 230.505 41.855 247.735 41.995 ;
		LAYER M4 ;
		RECT 71.735 38.390 88.965 40.270 ;
		LAYER M4 ;
		RECT 230.505 38.390 247.735 40.270 ;
		LAYER M4 ;
		RECT 548.045 45.460 565.275 47.505 ;
		LAYER M4 ;
		RECT 406.505 43.785 548.045 44.280 ;
		LAYER M4 ;
		RECT 0.000 47.415 654.735 53.235 ;
		LAYER M4 ;
		RECT 0.000 56.835 654.735 62.315 ;
		LAYER M4 ;
		RECT 247.735 34.505 389.275 35.000 ;
		LAYER M4 ;
		RECT 0.000 68.725 654.735 69.805 ;
		LAYER M4 ;
		RECT 0.000 78.005 654.345 79.085 ;
		LAYER M4 ;
		RECT 0.000 87.285 654.345 88.365 ;
		LAYER M4 ;
		RECT 0.000 42.325 654.735 43.405 ;
		LAYER M4 ;
		RECT 0.000 33.045 654.345 34.125 ;
		LAYER M4 ;
		RECT 0.000 96.565 654.345 97.645 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 654.555 102.850 ;
		LAYER M3 ;
		RECT 0.000 0.000 654.555 102.850 ;
		LAYER M2 ;
		RECT 0.000 0.000 654.555 102.850 ;
		LAYER M1 ;
		RECT 0.000 0.000 654.555 102.850 ;
		LAYER M2 ;
		RECT 654.555 54.680 654.735 54.760 ;
		LAYER VIA3 ;
		RECT 654.555 54.680 654.735 54.760 ;
		LAYER M1 ;
		RECT 654.555 46.460 654.735 46.580 ;
		LAYER VIA3 ;
		RECT 654.555 53.020 654.735 54.370 ;
		LAYER M1 ;
		RECT 654.555 54.660 654.735 54.780 ;
		LAYER M1 ;
		RECT 654.555 53.000 654.735 54.390 ;
		LAYER M3 ;
		RECT 654.555 50.970 654.735 52.320 ;
		LAYER M1 ;
		RECT 654.555 48.900 654.735 50.290 ;
		LAYER VIA3 ;
		RECT 654.555 48.530 654.735 48.610 ;
		LAYER VIA3 ;
		RECT 654.555 50.970 654.735 52.320 ;
		LAYER M1 ;
		RECT 654.555 50.560 654.735 50.680 ;
		LAYER VIA3 ;
		RECT 654.555 50.580 654.735 50.660 ;
		LAYER M1 ;
		RECT 654.555 46.850 654.735 48.240 ;
		LAYER M3 ;
		RECT 654.555 46.870 654.735 48.220 ;
		LAYER VIA3 ;
		RECT 654.555 46.870 654.735 48.220 ;
		LAYER M3 ;
		RECT 654.555 48.530 654.735 48.610 ;
		LAYER M1 ;
		RECT 654.555 44.950 654.735 46.190 ;
		LAYER M2 ;
		RECT 654.555 44.970 654.735 46.170 ;
		LAYER M3 ;
		RECT 654.555 44.970 654.735 46.170 ;
		LAYER VIA3 ;
		RECT 654.555 44.970 654.735 46.170 ;
		LAYER M2 ;
		RECT 654.555 46.480 654.735 46.560 ;
		LAYER M3 ;
		RECT 654.555 46.480 654.735 46.560 ;
		LAYER VIA3 ;
		RECT 654.555 46.480 654.735 46.560 ;
		LAYER VIA3 ;
		RECT 654.555 17.155 654.735 25.115 ;
		LAYER M1 ;
		RECT 654.555 17.135 654.735 25.135 ;
		LAYER M2 ;
		RECT 654.555 16.145 654.735 16.845 ;
		LAYER M1 ;
		RECT 654.555 16.125 654.735 16.865 ;
		LAYER M3 ;
		RECT 654.555 16.145 654.735 16.845 ;
		LAYER VIA3 ;
		RECT 654.555 16.145 654.735 16.845 ;
		LAYER M3 ;
		RECT 654.555 59.170 654.735 60.520 ;
		LAYER VIA3 ;
		RECT 654.555 57.120 654.735 58.470 ;
		LAYER M3 ;
		RECT 654.555 57.120 654.735 58.470 ;
		LAYER VIA3 ;
		RECT 654.555 59.170 654.735 60.520 ;
		LAYER M1 ;
		RECT 654.555 57.100 654.735 58.490 ;
		LAYER M1 ;
		RECT 654.555 44.235 654.735 44.680 ;
		LAYER VIA3 ;
		RECT 654.555 52.630 654.735 52.710 ;
		LAYER M2 ;
		RECT 654.555 48.530 654.735 48.610 ;
		LAYER M1 ;
		RECT 654.555 48.510 654.735 48.630 ;
		LAYER M2 ;
		RECT 654.555 46.870 654.735 48.220 ;
		LAYER M3 ;
		RECT 654.555 58.780 654.735 58.860 ;
		LAYER VIA3 ;
		RECT 654.555 58.780 654.735 58.860 ;
		LAYER M2 ;
		RECT 654.555 58.780 654.735 58.860 ;
		LAYER M1 ;
		RECT 654.555 58.760 654.735 58.880 ;
		LAYER M1 ;
		RECT 654.555 40.335 654.735 43.965 ;
		LAYER M2 ;
		RECT 654.555 40.355 654.735 43.945 ;
		LAYER VIA3 ;
		RECT 654.555 34.705 654.735 35.405 ;
		LAYER M3 ;
		RECT 654.555 54.680 654.735 54.760 ;
		LAYER M2 ;
		RECT 654.555 7.875 654.735 15.835 ;
		LAYER M1 ;
		RECT 654.555 7.855 654.735 15.855 ;
		LAYER M3 ;
		RECT 654.555 6.865 654.735 7.565 ;
		LAYER M2 ;
		RECT 654.555 6.865 654.735 7.565 ;
		LAYER M1 ;
		RECT 654.555 6.845 654.735 7.585 ;
		LAYER VIA3 ;
		RECT 654.555 6.865 654.735 7.565 ;
		LAYER M3 ;
		RECT 654.555 7.875 654.735 15.835 ;
		LAYER VIA3 ;
		RECT 654.555 7.875 654.735 15.835 ;
		LAYER M3 ;
		RECT 654.555 0.000 654.735 6.555 ;
		LAYER VIA3 ;
		RECT 654.555 0.000 654.735 6.555 ;
		LAYER M2 ;
		RECT 654.555 0.000 654.735 6.555 ;
		LAYER M1 ;
		RECT 654.555 0.000 654.735 6.575 ;
		LAYER VIA3 ;
		RECT 654.555 26.435 654.735 34.395 ;
		LAYER M2 ;
		RECT 654.555 34.705 654.735 35.405 ;
		LAYER M3 ;
		RECT 654.555 35.715 654.735 39.035 ;
		LAYER VIA3 ;
		RECT 654.555 35.715 654.735 39.035 ;
		LAYER M1 ;
		RECT 654.555 34.685 654.735 35.425 ;
		LAYER M1 ;
		RECT 654.555 35.695 654.735 39.055 ;
		LAYER M3 ;
		RECT 654.555 40.355 654.735 43.945 ;
		LAYER VIA3 ;
		RECT 654.555 40.355 654.735 43.945 ;
		LAYER VIA3 ;
		RECT 654.555 39.345 654.735 40.045 ;
		LAYER M3 ;
		RECT 654.555 39.345 654.735 40.045 ;
		LAYER M2 ;
		RECT 654.555 25.425 654.735 26.125 ;
		LAYER M3 ;
		RECT 654.555 25.425 654.735 26.125 ;
		LAYER M1 ;
		RECT 654.555 25.405 654.735 26.145 ;
		LAYER M3 ;
		RECT 654.555 17.155 654.735 25.115 ;
		LAYER VIA3 ;
		RECT 654.555 25.425 654.735 26.125 ;
		LAYER M2 ;
		RECT 654.555 17.155 654.735 25.115 ;
		LAYER M2 ;
		RECT 654.555 50.970 654.735 52.320 ;
		LAYER M2 ;
		RECT 654.555 48.920 654.735 50.270 ;
		LAYER M3 ;
		RECT 654.555 48.920 654.735 50.270 ;
		LAYER VIA3 ;
		RECT 654.555 48.920 654.735 50.270 ;
		LAYER M2 ;
		RECT 654.555 56.730 654.735 56.810 ;
		LAYER M3 ;
		RECT 654.555 56.730 654.735 56.810 ;
		LAYER M1 ;
		RECT 654.555 55.050 654.735 56.440 ;
		LAYER VIA3 ;
		RECT 654.555 56.730 654.735 56.810 ;
		LAYER VIA3 ;
		RECT 654.555 55.070 654.735 56.420 ;
		LAYER M2 ;
		RECT 654.555 44.255 654.735 44.660 ;
		LAYER M3 ;
		RECT 654.555 44.255 654.735 44.660 ;
		LAYER VIA3 ;
		RECT 654.555 44.255 654.735 44.660 ;
		LAYER M4 ;
		RECT 389.275 98.025 406.505 98.555 ;
		LAYER M4 ;
		RECT 389.275 99.700 406.505 101.745 ;
		LAYER M4 ;
		RECT 389.275 71.860 406.505 73.905 ;
		LAYER M4 ;
		RECT 389.275 68.255 406.505 68.395 ;
		LAYER M4 ;
		RECT 389.275 64.790 406.505 66.670 ;
		LAYER M4 ;
		RECT 389.275 83.350 406.505 85.230 ;
		LAYER M4 ;
		RECT 389.275 81.140 406.505 83.185 ;
		LAYER M4 ;
		RECT 389.275 70.185 406.505 70.715 ;
		LAYER M4 ;
		RECT 389.275 96.095 406.505 96.235 ;
		LAYER M4 ;
		RECT 389.275 77.535 406.505 77.675 ;
		LAYER M4 ;
		RECT 389.275 74.070 406.505 75.950 ;
		LAYER M4 ;
		RECT 389.275 92.630 406.505 94.510 ;
		LAYER M4 ;
		RECT 389.275 86.815 406.505 86.955 ;
		LAYER M4 ;
		RECT 389.275 88.745 406.505 89.275 ;
		LAYER M4 ;
		RECT 389.275 90.420 406.505 92.465 ;
		LAYER M4 ;
		RECT 389.275 79.465 406.505 79.995 ;
		LAYER M4 ;
		RECT 71.735 29.110 88.965 30.990 ;
		LAYER M4 ;
		RECT 71.735 26.900 88.965 28.945 ;
		LAYER M4 ;
		RECT 71.735 25.225 88.965 25.755 ;
		LAYER M4 ;
		RECT 71.735 19.830 88.965 21.710 ;
		LAYER M4 ;
		RECT 71.735 23.295 88.965 23.435 ;
		LAYER M4 ;
		RECT 71.735 32.575 88.965 32.715 ;
		LAYER M4 ;
		RECT 71.735 17.620 88.965 19.665 ;
		LAYER M4 ;
		RECT 71.735 10.550 88.965 12.430 ;
		LAYER M4 ;
		RECT 71.735 14.015 88.965 14.155 ;
		LAYER M4 ;
		RECT 71.735 15.945 88.965 16.475 ;
		LAYER M4 ;
		RECT 389.275 15.945 406.505 16.475 ;
		LAYER M4 ;
		RECT 389.275 17.620 406.505 19.665 ;
		LAYER M4 ;
		RECT 230.505 32.575 247.735 32.715 ;
		LAYER M4 ;
		RECT 389.275 32.575 406.505 32.715 ;
		LAYER M4 ;
		RECT 247.735 25.225 389.275 25.720 ;
		LAYER M4 ;
		RECT 389.275 10.550 406.505 12.430 ;
		LAYER M4 ;
		RECT 88.965 15.945 230.505 16.440 ;
		LAYER M4 ;
		RECT 230.505 15.945 247.735 16.475 ;
		LAYER M4 ;
		RECT 230.505 17.620 247.735 19.665 ;
		LAYER M4 ;
		RECT 230.505 10.550 247.735 12.430 ;
		LAYER M4 ;
		RECT 230.505 14.015 247.735 14.155 ;
		LAYER M4 ;
		RECT 88.965 25.225 230.505 25.720 ;
		LAYER M4 ;
		RECT 230.505 25.225 247.735 25.755 ;
		LAYER M4 ;
		RECT 230.505 23.295 247.735 23.435 ;
		LAYER M4 ;
		RECT 230.505 19.830 247.735 21.710 ;
		LAYER M4 ;
		RECT 230.505 29.110 247.735 30.990 ;
		LAYER M4 ;
		RECT 230.505 26.900 247.735 28.945 ;
		LAYER M4 ;
		RECT 0.000 14.015 1.365 14.155 ;
		LAYER M4 ;
		RECT 0.000 23.295 1.365 23.435 ;
		LAYER M4 ;
		RECT 0.000 25.225 71.735 25.720 ;
		LAYER M4 ;
		RECT 0.000 15.945 71.735 16.440 ;
		LAYER M4 ;
		RECT 88.965 34.505 230.505 35.000 ;
		LAYER M4 ;
		RECT 230.505 34.505 247.735 35.035 ;
		LAYER M4 ;
		RECT 230.505 36.180 247.735 38.225 ;
		LAYER M4 ;
		RECT 389.275 38.390 406.505 40.270 ;
		LAYER M4 ;
		RECT 389.275 41.855 406.505 41.995 ;
		LAYER M4 ;
		RECT 389.275 43.785 406.505 44.315 ;
		LAYER M4 ;
		RECT 389.275 45.460 406.505 47.505 ;
		LAYER M4 ;
		RECT 247.735 88.745 389.275 89.240 ;
		LAYER M4 ;
		RECT 247.735 98.025 389.275 98.520 ;
		LAYER M4 ;
		RECT 247.735 79.465 389.275 79.960 ;
		LAYER M4 ;
		RECT 247.735 70.185 389.275 70.680 ;
		LAYER M4 ;
		RECT 0.000 77.535 1.365 77.675 ;
		LAYER M4 ;
		RECT 0.000 79.465 71.735 79.960 ;
		LAYER M4 ;
		RECT 0.000 70.185 71.735 70.680 ;
		LAYER M4 ;
		RECT 0.000 86.815 1.365 86.955 ;
		LAYER M4 ;
		RECT 0.000 96.095 1.365 96.235 ;
		LAYER M4 ;
		RECT 0.000 88.745 71.735 89.240 ;
		LAYER M4 ;
		RECT 0.000 98.025 71.735 98.520 ;
		LAYER M4 ;
		RECT 71.735 98.025 88.965 98.555 ;
		LAYER M4 ;
		RECT 71.735 96.095 88.965 96.235 ;
		LAYER M4 ;
		RECT 71.735 92.630 88.965 94.510 ;
		LAYER M4 ;
		RECT 71.735 90.420 88.965 92.465 ;
		LAYER M4 ;
		RECT 71.735 99.700 88.965 101.745 ;
		LAYER M4 ;
		RECT 71.735 83.350 88.965 85.230 ;
		LAYER M4 ;
		RECT 71.735 86.815 88.965 86.955 ;
		LAYER M4 ;
		RECT 71.735 88.745 88.965 89.275 ;
		LAYER M4 ;
		RECT 230.505 99.700 247.735 101.745 ;
		LAYER M4 ;
		RECT 230.505 88.745 247.735 89.275 ;
		LAYER M4 ;
		RECT 230.505 86.815 247.735 86.955 ;
		LAYER M4 ;
		RECT 230.505 83.350 247.735 85.230 ;
		LAYER M4 ;
		RECT 230.505 81.140 247.735 83.185 ;
		LAYER M4 ;
		RECT 230.505 74.070 247.735 75.950 ;
		LAYER M4 ;
		RECT 230.505 77.535 247.735 77.675 ;
		LAYER M4 ;
		RECT 230.505 71.860 247.735 73.905 ;
		LAYER M4 ;
		RECT 230.505 70.185 247.735 70.715 ;
		LAYER M4 ;
		RECT 71.735 79.465 88.965 79.995 ;
		LAYER M4 ;
		RECT 71.735 81.140 88.965 83.185 ;
		LAYER M4 ;
		RECT 88.965 98.025 230.505 98.520 ;
		LAYER M4 ;
		RECT 88.965 88.745 230.505 89.240 ;
		LAYER M4 ;
		RECT 71.735 77.535 88.965 77.675 ;
		LAYER M4 ;
		RECT 71.735 74.070 88.965 75.950 ;
		LAYER M4 ;
		RECT 71.735 71.860 88.965 73.905 ;
		LAYER M4 ;
		RECT 71.735 70.185 88.965 70.715 ;
		LAYER M4 ;
		RECT 230.505 98.025 247.735 98.555 ;
		LAYER M4 ;
		RECT 230.505 96.095 247.735 96.235 ;
		LAYER M4 ;
		RECT 230.505 92.630 247.735 94.510 ;
		LAYER M4 ;
		RECT 230.505 90.420 247.735 92.465 ;
		LAYER M4 ;
		RECT 88.965 79.465 230.505 79.960 ;
		LAYER M4 ;
		RECT 230.505 79.465 247.735 79.995 ;
		LAYER M4 ;
		RECT 88.965 70.185 230.505 70.680 ;
		LAYER M4 ;
		RECT 318.855 63.465 353.415 64.420 ;
		LAYER M4 ;
		RECT 318.155 62.885 318.855 64.420 ;
		LAYER M4 ;
		RECT 283.595 63.465 318.155 64.420 ;
		LAYER M4 ;
		RECT 248.875 63.465 282.895 64.420 ;
		LAYER M4 ;
		RECT 230.505 64.790 247.735 66.670 ;
		LAYER M4 ;
		RECT 230.505 68.255 247.735 68.395 ;
		LAYER M4 ;
		RECT 248.335 62.885 318.155 63.465 ;
		LAYER M4 ;
		RECT 229.905 62.885 248.335 64.420 ;
		LAYER M4 ;
		RECT 89.565 62.885 159.385 63.465 ;
		LAYER M4 ;
		RECT 160.085 62.885 229.905 63.465 ;
		LAYER M4 ;
		RECT 195.345 63.465 229.905 64.420 ;
		LAYER M4 ;
		RECT 160.085 63.465 194.645 64.420 ;
		LAYER M4 ;
		RECT 159.385 62.885 160.085 64.420 ;
		LAYER M4 ;
		RECT 124.825 63.465 159.385 64.420 ;
		LAYER M4 ;
		RECT 71.735 64.790 88.965 66.670 ;
		LAYER M4 ;
		RECT 71.735 68.255 88.965 68.395 ;
		LAYER M4 ;
		RECT 90.105 63.465 124.125 64.420 ;
		LAYER M4 ;
		RECT 1.315 63.465 35.875 64.420 ;
		LAYER M4 ;
		RECT 36.575 63.465 71.135 64.420 ;
		LAYER M4 ;
		RECT 1.315 62.885 71.135 63.465 ;
		LAYER M4 ;
		RECT 71.135 62.885 89.565 64.420 ;
		LAYER M4 ;
		RECT 0.000 62.885 1.315 64.420 ;
		LAYER M4 ;
		RECT 0.000 68.255 1.365 68.395 ;
		LAYER M4 ;
		RECT 0.000 32.575 1.365 32.715 ;
		LAYER M4 ;
		RECT 0.000 41.855 1.365 41.995 ;
		LAYER M4 ;
		RECT 0.000 43.785 71.735 44.280 ;
		LAYER M4 ;
		RECT 71.735 36.180 88.965 38.225 ;
		LAYER M4 ;
		RECT 71.735 34.505 88.965 35.035 ;
		LAYER M4 ;
		RECT 0.000 34.505 71.735 35.000 ;
		LAYER M4 ;
		RECT 354.115 63.465 374.095 64.420 ;
		LAYER M4 ;
		RECT 318.855 62.885 374.095 63.465 ;
		LAYER M4 ;
		RECT 247.735 43.785 389.275 44.280 ;
		LAYER M4 ;
		RECT 71.735 43.785 88.965 44.315 ;
		LAYER M4 ;
		RECT 71.735 45.460 88.965 47.505 ;
		LAYER M4 ;
		RECT 230.505 43.785 247.735 44.315 ;
		LAYER M4 ;
		RECT 230.505 45.460 247.735 47.505 ;
		LAYER M4 ;
		RECT 88.965 43.785 230.505 44.280 ;
	END
	# End of OBS

END TS1N28HPCPHVTB32768X9M16SSO

END LIBRARY
