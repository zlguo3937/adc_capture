// Copyright (c) 2024 by JLSemi Inc.
// --------------------------------------------------------------------
//
//                     JLSemi
//                     Shanghai, China
//                     Name : Zhiling Guo
//                     Email: zlguo@jlsemi.com
//
// --------------------------------------------------------------------
// --------------------------------------------------------------------
//  Revision History:1.0
//  Date          By            Revision    Design Description
//---------------------------------------------------------------------
//  2024-05-06    zlguo         1.0         package_gen
// --------------------------------------------------------------------
// --------------------------------------------------------------------
module package_gen
(
    output  wire    [35:0]  pkt_gen_data_0,
    output  wire    [35:0]  pkt_gen_data_1,
    output  wire    [35:0]  pkt_gen_data_2,
    output  wire    [35:0]  pkt_gen_data_3,
    output  wire    [35:0]  pkt_gen_data_4,
    output  wire    [35:0]  pkt_gen_data_5,
    output  wire    [35:0]  pkt_gen_data_6,
    output  wire    [35:0]  pkt_gen_data_7,
    output  wire    [35:0]  pkt_gen_data_8,
    output  wire    [35:0]  pkt_gen_data_9,
    output  wire    [35:0]  pkt_gen_data_10,
    output  wire    [35:0]  pkt_gen_data_11,
    output  wire    [35:0]  pkt_gen_data_12,
    output  wire    [35:0]  pkt_gen_data_13,
    output  wire    [35:0]  pkt_gen_data_14,
    output  wire    [35:0]  pkt_gen_data_15,
    output  wire    [35:0]  pkt_gen_data_16,
    output  wire    [35:0]  pkt_gen_data_17,
    output  wire    [35:0]  pkt_gen_data_18,
    output  wire    [35:0]  pkt_gen_data_19,
    output  wire    [35:0]  pkt_gen_data_20,
    output  wire    [35:0]  pkt_gen_data_21,
    output  wire    [35:0]  pkt_gen_data_22,
    output  wire    [35:0]  pkt_gen_data_23,

    output  wire    [35:0]  pkt_gen_48data_0,
    output  wire    [35:0]  pkt_gen_48data_1,
    output  wire    [35:0]  pkt_gen_48data_2,
    output  wire    [35:0]  pkt_gen_48data_3,
    output  wire    [35:0]  pkt_gen_48data_4,
    output  wire    [35:0]  pkt_gen_48data_5,
    output  wire    [35:0]  pkt_gen_48data_6,
    output  wire    [35:0]  pkt_gen_48data_7,
    output  wire    [35:0]  pkt_gen_48data_8,
    output  wire    [35:0]  pkt_gen_48data_9,
    output  wire    [35:0]  pkt_gen_48data_10,
    output  wire    [35:0]  pkt_gen_48data_11

);

endmodule
