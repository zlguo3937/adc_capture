// Copyright (c) 2024 by JLSemi Inc.
// --------------------------------------------------------------------
//
//                     JLSemi
//                     Shanghai, China
//                     Name : Zhiling Guo
//                     Email: zlguo@jlsemi.com
//
// --------------------------------------------------------------------
// --------------------------------------------------------------------
//  Revision History:1.0
//  Date          By            Revision    Design Description
//---------------------------------------------------------------------
//  2024-05-06    zlguo         1.0         DIGITAL_WRAPPER
// --------------------------------------------------------------------
// --------------------------------------------------------------------
`timescale 1ns/1ns
module DIGITAL_WRAPPER
(
    input   wire            CLK200M,
    input   wire            ADC_CLK500M,
    input   wire            ADC48_CLK500M,

    input   wire    [8:0]   ADC_DATA_0 ,
    input   wire    [8:0]   ADC_DATA_1 ,
    input   wire    [8:0]   ADC_DATA_2 ,
    input   wire    [8:0]   ADC_DATA_3 ,
    input   wire    [8:0]   ADC_DATA_4 ,
    input   wire    [8:0]   ADC_DATA_5 ,
    input   wire    [8:0]   ADC_DATA_6 ,
    input   wire    [8:0]   ADC_DATA_7 ,
    input   wire    [8:0]   ADC_DATA_8 ,
    input   wire    [8:0]   ADC_DATA_9 ,
    input   wire    [8:0]   ADC_DATA_10,
    input   wire    [8:0]   ADC_DATA_11,
    input   wire    [8:0]   ADC_DATA_12,
    input   wire    [8:0]   ADC_DATA_13,
    input   wire    [8:0]   ADC_DATA_14,
    input   wire    [8:0]   ADC_DATA_15,
    input   wire    [8:0]   ADC_DATA_16,
    input   wire    [8:0]   ADC_DATA_17,
    input   wire    [8:0]   ADC_DATA_18,
    input   wire    [8:0]   ADC_DATA_19,
    input   wire    [8:0]   ADC_DATA_20,
    input   wire    [8:0]   ADC_DATA_21,
    input   wire    [8:0]   ADC_DATA_22,
    input   wire    [8:0]   ADC_DATA_23,
    input   wire    [8:0]   ADC_DATA_24,
    input   wire    [8:0]   ADC_DATA_25,
    input   wire    [8:0]   ADC_DATA_26,
    input   wire    [8:0]   ADC_DATA_27,
    input   wire    [8:0]   ADC_DATA_28,
    input   wire    [8:0]   ADC_DATA_29,
    input   wire    [8:0]   ADC_DATA_30,
    input   wire    [8:0]   ADC_DATA_31,
    input   wire    [8:0]   ADC_DATA_32,
    input   wire    [8:0]   ADC_DATA_33,
    input   wire    [8:0]   ADC_DATA_34,
    input   wire    [8:0]   ADC_DATA_35,
    input   wire    [8:0]   ADC_DATA_36,
    input   wire    [8:0]   ADC_DATA_37,
    input   wire    [8:0]   ADC_DATA_38,
    input   wire    [8:0]   ADC_DATA_39,
    input   wire    [8:0]   ADC_DATA_40,
    input   wire    [8:0]   ADC_DATA_41,
    input   wire    [8:0]   ADC_DATA_42,
    input   wire    [8:0]   ADC_DATA_43,
    input   wire    [8:0]   ADC_DATA_44,
    input   wire    [8:0]   ADC_DATA_45,
    input   wire    [8:0]   ADC_DATA_46,
    input   wire    [8:0]   ADC_DATA_47,
    input   wire    [8:0]   ADC_DATA_48,
    input   wire    [8:0]   ADC_DATA_49,
    input   wire    [8:0]   ADC_DATA_50,
    input   wire    [8:0]   ADC_DATA_51,
    input   wire    [8:0]   ADC_DATA_52,
    input   wire    [8:0]   ADC_DATA_53,
    input   wire    [8:0]   ADC_DATA_54,
    input   wire    [8:0]   ADC_DATA_55,
    input   wire    [8:0]   ADC_DATA_56,
    input   wire    [8:0]   ADC_DATA_57,
    input   wire    [8:0]   ADC_DATA_58,
    input   wire    [8:0]   ADC_DATA_59,
    input   wire    [8:0]   ADC_DATA_60,
    input   wire    [8:0]   ADC_DATA_61,
    input   wire    [8:0]   ADC_DATA_62,
    input   wire    [8:0]   ADC_DATA_63,
    input   wire    [8:0]   ADC_DATA_64,
    input   wire    [8:0]   ADC_DATA_65,
    input   wire    [8:0]   ADC_DATA_66,
    input   wire    [8:0]   ADC_DATA_67,
    input   wire    [8:0]   ADC_DATA_68,
    input   wire    [8:0]   ADC_DATA_69,
    input   wire    [8:0]   ADC_DATA_70,
    input   wire    [8:0]   ADC_DATA_71,
    input   wire    [8:0]   ADC_DATA_72,
    input   wire    [8:0]   ADC_DATA_73,
    input   wire    [8:0]   ADC_DATA_74,
    input   wire    [8:0]   ADC_DATA_75,
    input   wire    [8:0]   ADC_DATA_76,
    input   wire    [8:0]   ADC_DATA_77,
    input   wire    [8:0]   ADC_DATA_78,
    input   wire    [8:0]   ADC_DATA_79,
    input   wire    [8:0]   ADC_DATA_80,
    input   wire    [8:0]   ADC_DATA_81,
    input   wire    [8:0]   ADC_DATA_82,
    input   wire    [8:0]   ADC_DATA_83,
    input   wire    [8:0]   ADC_DATA_84,
    input   wire    [8:0]   ADC_DATA_85,
    input   wire    [8:0]   ADC_DATA_86,
    input   wire    [8:0]   ADC_DATA_87,
    input   wire    [8:0]   ADC_DATA_88,
    input   wire    [8:0]   ADC_DATA_89,
    input   wire    [8:0]   ADC_DATA_90,
    input   wire    [8:0]   ADC_DATA_91,
    input   wire    [8:0]   ADC_DATA_92,
    input   wire    [8:0]   ADC_DATA_93,
    input   wire    [8:0]   ADC_DATA_94,
    input   wire    [8:0]   ADC_DATA_95,
    input   wire    [8:0]   ADC48_DATA_0,
    input   wire    [8:0]   ADC48_DATA_1,
    input   wire    [8:0]   ADC48_DATA_2,
    input   wire    [8:0]   ADC48_DATA_3,
    input   wire    [8:0]   ADC48_DATA_4,
    input   wire    [8:0]   ADC48_DATA_5,
    input   wire    [8:0]   ADC48_DATA_6,
    input   wire    [8:0]   ADC48_DATA_7,
    input   wire    [8:0]   ADC48_DATA_8,
    input   wire    [8:0]   ADC48_DATA_9,
    input   wire    [8:0]   ADC48_DATA_10,
    input   wire    [8:0]   ADC48_DATA_11,
    input   wire    [8:0]   ADC48_DATA_12,
    input   wire    [8:0]   ADC48_DATA_13,
    input   wire    [8:0]   ADC48_DATA_14,
    input   wire    [8:0]   ADC48_DATA_15,
    input   wire    [8:0]   ADC48_DATA_16,
    input   wire    [8:0]   ADC48_DATA_17,
    input   wire    [8:0]   ADC48_DATA_18,
    input   wire    [8:0]   ADC48_DATA_19,
    input   wire    [8:0]   ADC48_DATA_20,
    input   wire    [8:0]   ADC48_DATA_21,
    input   wire    [8:0]   ADC48_DATA_22,
    input   wire    [8:0]   ADC48_DATA_23,
    input   wire    [8:0]   ADC48_DATA_24,
    input   wire    [8:0]   ADC48_DATA_25,
    input   wire    [8:0]   ADC48_DATA_26,
    input   wire    [8:0]   ADC48_DATA_27,
    input   wire    [8:0]   ADC48_DATA_28,
    input   wire    [8:0]   ADC48_DATA_29,
    input   wire    [8:0]   ADC48_DATA_30,
    input   wire    [8:0]   ADC48_DATA_31,
    input   wire    [8:0]   ADC48_DATA_32,
    input   wire    [8:0]   ADC48_DATA_33,
    input   wire    [8:0]   ADC48_DATA_34,
    input   wire    [8:0]   ADC48_DATA_35,
    input   wire    [8:0]   ADC48_DATA_36,
    input   wire    [8:0]   ADC48_DATA_37,
    input   wire    [8:0]   ADC48_DATA_38,
    input   wire    [8:0]   ADC48_DATA_39,
    input   wire    [8:0]   ADC48_DATA_40,
    input   wire    [8:0]   ADC48_DATA_41,
    input   wire    [8:0]   ADC48_DATA_42,
    input   wire    [8:0]   ADC48_DATA_43,
    input   wire    [8:0]   ADC48_DATA_44,
    input   wire    [8:0]   ADC48_DATA_45,
    input   wire    [8:0]   ADC48_DATA_46,
    input   wire    [8:0]   ADC48_DATA_47,

    inout   wire            PAD1_ADC_DATA_1,
    inout   wire            PAD2_ADC_DATA_2,
    inout   wire            PAD3_ADC_DATA_3,
    inout   wire            PAD4_ADC_DATA_4,
    inout   wire            PAD5_ADC_DATA_5,
    inout   wire            PAD6_ADC_DATA_6,
    inout   wire            PAD7_ADC_DATA_7,
    inout   wire            PAD8_ADC_DATA_8,
    inout   wire            PAD9_ADC_DATA_9,
    inout   wire            PAD10_ADC_DATA_10,
    inout   wire            PAD11_ADC_DATA_11,
    inout   wire            PAD12_ADC_DATA_12,
    inout   wire            PAD13_ADC_DATA_13,
    inout   wire            PAD14_ADC_DATA_14,
    inout   wire            PAD15_ADC_DATA_15,
    inout   wire            PAD16_ADC_DATA_16,
    inout   wire            PAD17_ADC_DATA_17,
    inout   wire            PAD18_ADC_DATA_18,
    inout   wire            PAD19_ADC_DATA_VALID,
    inout   wire            PAD20_RSTN,
    inout   wire            PAD21_CLK_RD,
    inout   wire            PAD22_MDC,
    inout   wire            PAD23_MDIO
);

    // analog_signal_mux
    wire            ANA_CLK200M;
    wire            ANA_ADC_CLK500M;
    wire            ANA_ADC48_CLK500M;
    wire    [35:0]  ANA_ADC_DATA_0;
    wire    [35:0]  ANA_ADC_DATA_1;
    wire    [35:0]  ANA_ADC_DATA_2;
    wire    [35:0]  ANA_ADC_DATA_3;
    wire    [35:0]  ANA_ADC_DATA_4;
    wire    [35:0]  ANA_ADC_DATA_5;
    wire    [35:0]  ANA_ADC_DATA_6;
    wire    [35:0]  ANA_ADC_DATA_7;
    wire    [35:0]  ANA_ADC_DATA_8;
    wire    [35:0]  ANA_ADC_DATA_9;
    wire    [35:0]  ANA_ADC_DATA_10;
    wire    [35:0]  ANA_ADC_DATA_11;
    wire    [35:0]  ANA_ADC_DATA_12;
    wire    [35:0]  ANA_ADC_DATA_13;
    wire    [35:0]  ANA_ADC_DATA_14;
    wire    [35:0]  ANA_ADC_DATA_15;
    wire    [35:0]  ANA_ADC_DATA_16;
    wire    [35:0]  ANA_ADC_DATA_17;
    wire    [35:0]  ANA_ADC_DATA_18;
    wire    [35:0]  ANA_ADC_DATA_19;
    wire    [35:0]  ANA_ADC_DATA_20;
    wire    [35:0]  ANA_ADC_DATA_21;
    wire    [35:0]  ANA_ADC_DATA_22;
    wire    [35:0]  ANA_ADC_DATA_23;

    wire    [35:0]  ANA_ADC48_DATA_0;
    wire    [35:0]  ANA_ADC48_DATA_1;
    wire    [35:0]  ANA_ADC48_DATA_2;
    wire    [35:0]  ANA_ADC48_DATA_3;
    wire    [35:0]  ANA_ADC48_DATA_4;
    wire    [35:0]  ANA_ADC48_DATA_5;
    wire    [35:0]  ANA_ADC48_DATA_6;
    wire    [35:0]  ANA_ADC48_DATA_7;
    wire    [35:0]  ANA_ADC48_DATA_8;
    wire    [35:0]  ANA_ADC48_DATA_9;
    wire    [35:0]  ANA_ADC48_DATA_10;
    wire    [35:0]  ANA_ADC48_DATA_11;

    // crg
    wire    [8:0]   rf_pktctrl_gap;
    wire    [8:0]   rf_pktctrl_phase;
    wire            rf_pktctrl_clk_en;
    wire            rf_pktctrl_sw_rstn;
    wire            pktctrl_clk;
    wire            pktctrl_rstn;
    wire            clk_200m;
    wire            rstn_200m;
    wire            adc96_rstn;
    wire            adc48_rstn;

    // io pad
    wire            CLK_RD;
    wire            DATA_RD_EN; 
    wire            RSTN; 

    wire    [17:0]  ADC_DATA;
    wire            ADC_DATA_VALID;
    wire            MDIO;
    wire            MDC;
    wire            mdio_out;
    wire            mdio_oen;

    // ctrl_sys
    wire            rf_self_test_mode;

    wire            rf_capture_mode;
    wire            rf_capture_start;
    wire            rf_capture_again;

    wire            rf_96path_en;
    wire    [1:0]   rf_pkt_data_length;
    wire    [15:0]  rf_pkt_idle_length;

    wire    [6:0]   rf_mdio_data_sel;
    wire    [14:0]  rf_mdio_memory_addr;
    wire    [8:0]   rf_mdio_pkt_data;

    wire            tri_succeed     ;
    wire    [31:0]  tri_data        ;
    wire            tri_data_vld    ;

    wire            capture_enable  ;
    wire            capture_start   ;

    wire    [3:0]   capture_mode    ;
    wire    [12:0]  capture_max_addr;
    wire    [12:0]  pre_trigger_num ;

    wire    [15:0]  trigger_pattern0;
    wire    [15:0]  trigger_pattern1;
    wire    [15:0]  trigger_mode0   ;
    wire    [15:0]  trigger_mode1   ;
    wire    [15:0]  trigger_mode2   ;
    wire    [15:0]  trigger_mode3   ;
    wire    [15:0]  trigger_mode4   ;
    wire    [15:0]  trigger_mode5   ;
    wire    [15:0]  trigger_logic0  ;
    wire    [15:0]  trigger_logic1  ;
    wire            store_mode      ;

    wire    [12:0]  read_start_addr ;
    wire    [12:0]  tri_addr        ;
    wire            capture_done_rd ;
    wire            capture_done    ;

    wire            tri_succeed_cnt_overflow_mode;
    wire            tri_succeed_cnt_clr;
    wire    [7:0]   tri_succeed_cnt ;

    wire            capture_rd_en   ;
    wire    [12:0]  capture_rd_addr ;
    wire    [15:0]  capture_rd_data0;
    wire    [15:0]  capture_rd_data1;

    wire    [15:0]  write_info      ; // write_en + waddr --> 1bit + 15bit
    wire            write_done      ; // write_done

    wire    [12:0]  pkt_ctrl_info   ; // main_fsm: 1bit-write_en + 1bit-wr_done + 1bit-fast_read_en + 5bit-curr_sta + 5bit-next_sta
    wire    [15:0]  fast_info       ; // fast_read_en + fast_raddr --> 1bit + 15bit
    wire            fast_rd_done    ; // fast_rd_done

    wire    [13:0]  fast_main_fsm   ; // 7bit-curr_sta + 7bit-next_sta
    wire    [5:0]   fast_pkt_fsm    ; // pkt_en + read_en + 2bit-curr_sta + 2bit-next_sta
    wire    [15:0]  idle_cnt        ; // idle_cnt
    wire    [9:0]   RD_info         ; // RD + RD_CNT

    // analog_signal_mux instantiation
    analog_signal_mux
    u_analog_signal_mux
    (
    .adc96_rstn                 (adc96_rstn                 ),
    .adc48_rstn                 (adc48_rstn                 ),
    .CLK200M                    (CLK200M                    ),
    .ADC_CLK500M                (ADC_CLK500M                ),
    .ADC48_CLK500M              (ADC48_CLK500M              ),

    .ADC_DATA_0                 (ADC_DATA_0                 ),
    .ADC_DATA_1                 (ADC_DATA_1                 ),
    .ADC_DATA_2                 (ADC_DATA_2                 ),
    .ADC_DATA_3                 (ADC_DATA_3                 ),
    .ADC_DATA_4                 (ADC_DATA_4                 ),
    .ADC_DATA_5                 (ADC_DATA_5                 ),
    .ADC_DATA_6                 (ADC_DATA_6                 ),
    .ADC_DATA_7                 (ADC_DATA_7                 ),
    .ADC_DATA_8                 (ADC_DATA_8                 ),
    .ADC_DATA_9                 (ADC_DATA_9                 ),
    .ADC_DATA_10                (ADC_DATA_10                ),
    .ADC_DATA_11                (ADC_DATA_11                ),
    .ADC_DATA_12                (ADC_DATA_12                ),
    .ADC_DATA_13                (ADC_DATA_13                ),
    .ADC_DATA_14                (ADC_DATA_14                ),
    .ADC_DATA_15                (ADC_DATA_15                ),
    .ADC_DATA_16                (ADC_DATA_16                ),
    .ADC_DATA_17                (ADC_DATA_17                ),
    .ADC_DATA_18                (ADC_DATA_18                ),
    .ADC_DATA_19                (ADC_DATA_19                ),
    .ADC_DATA_20                (ADC_DATA_20                ),
    .ADC_DATA_21                (ADC_DATA_21                ),
    .ADC_DATA_22                (ADC_DATA_22                ),
    .ADC_DATA_23                (ADC_DATA_23                ),
    .ADC_DATA_24                (ADC_DATA_24                ),
    .ADC_DATA_25                (ADC_DATA_25                ),
    .ADC_DATA_26                (ADC_DATA_26                ),
    .ADC_DATA_27                (ADC_DATA_27                ),
    .ADC_DATA_28                (ADC_DATA_28                ),
    .ADC_DATA_29                (ADC_DATA_29                ),
    .ADC_DATA_30                (ADC_DATA_30                ),
    .ADC_DATA_31                (ADC_DATA_31                ),
    .ADC_DATA_32                (ADC_DATA_32                ),
    .ADC_DATA_33                (ADC_DATA_33                ),
    .ADC_DATA_34                (ADC_DATA_34                ),
    .ADC_DATA_35                (ADC_DATA_35                ),
    .ADC_DATA_36                (ADC_DATA_36                ),
    .ADC_DATA_37                (ADC_DATA_37                ),
    .ADC_DATA_38                (ADC_DATA_38                ),
    .ADC_DATA_39                (ADC_DATA_39                ),
    .ADC_DATA_40                (ADC_DATA_40                ),
    .ADC_DATA_41                (ADC_DATA_41                ),
    .ADC_DATA_42                (ADC_DATA_42                ),
    .ADC_DATA_43                (ADC_DATA_43                ),
    .ADC_DATA_44                (ADC_DATA_44                ),
    .ADC_DATA_45                (ADC_DATA_45                ),
    .ADC_DATA_46                (ADC_DATA_46                ),
    .ADC_DATA_47                (ADC_DATA_47                ),
    .ADC_DATA_48                (ADC_DATA_48                ),
    .ADC_DATA_49                (ADC_DATA_49                ),
    .ADC_DATA_50                (ADC_DATA_50                ),
    .ADC_DATA_51                (ADC_DATA_51                ),
    .ADC_DATA_52                (ADC_DATA_52                ),
    .ADC_DATA_53                (ADC_DATA_53                ),
    .ADC_DATA_54                (ADC_DATA_54                ),
    .ADC_DATA_55                (ADC_DATA_55                ),
    .ADC_DATA_56                (ADC_DATA_56                ),
    .ADC_DATA_57                (ADC_DATA_57                ),
    .ADC_DATA_58                (ADC_DATA_58                ),
    .ADC_DATA_59                (ADC_DATA_59                ),
    .ADC_DATA_60                (ADC_DATA_60                ),
    .ADC_DATA_61                (ADC_DATA_61                ),
    .ADC_DATA_62                (ADC_DATA_62                ),
    .ADC_DATA_63                (ADC_DATA_63                ),
    .ADC_DATA_64                (ADC_DATA_64                ),
    .ADC_DATA_65                (ADC_DATA_65                ),
    .ADC_DATA_66                (ADC_DATA_66                ),
    .ADC_DATA_67                (ADC_DATA_67                ),
    .ADC_DATA_68                (ADC_DATA_68                ),
    .ADC_DATA_69                (ADC_DATA_69                ),
    .ADC_DATA_70                (ADC_DATA_70                ),
    .ADC_DATA_71                (ADC_DATA_71                ),
    .ADC_DATA_72                (ADC_DATA_72                ),
    .ADC_DATA_73                (ADC_DATA_73                ),
    .ADC_DATA_74                (ADC_DATA_74                ),
    .ADC_DATA_75                (ADC_DATA_75                ),
    .ADC_DATA_76                (ADC_DATA_76                ),
    .ADC_DATA_77                (ADC_DATA_77                ),
    .ADC_DATA_78                (ADC_DATA_78                ),
    .ADC_DATA_79                (ADC_DATA_79                ),
    .ADC_DATA_80                (ADC_DATA_80                ),
    .ADC_DATA_81                (ADC_DATA_81                ),
    .ADC_DATA_82                (ADC_DATA_82                ),
    .ADC_DATA_83                (ADC_DATA_83                ),
    .ADC_DATA_84                (ADC_DATA_84                ),
    .ADC_DATA_85                (ADC_DATA_85                ),
    .ADC_DATA_86                (ADC_DATA_86                ),
    .ADC_DATA_87                (ADC_DATA_87                ),
    .ADC_DATA_88                (ADC_DATA_88                ),
    .ADC_DATA_89                (ADC_DATA_89                ),
    .ADC_DATA_90                (ADC_DATA_90                ),
    .ADC_DATA_91                (ADC_DATA_91                ),
    .ADC_DATA_92                (ADC_DATA_92                ),
    .ADC_DATA_93                (ADC_DATA_93                ),
    .ADC_DATA_94                (ADC_DATA_94                ),
    .ADC_DATA_95                (ADC_DATA_95                ),
    .ADC48_DATA_0               (ADC48_DATA_0               ),
    .ADC48_DATA_1               (ADC48_DATA_1               ),
    .ADC48_DATA_2               (ADC48_DATA_2               ),
    .ADC48_DATA_3               (ADC48_DATA_3               ),
    .ADC48_DATA_4               (ADC48_DATA_4               ),
    .ADC48_DATA_5               (ADC48_DATA_5               ),
    .ADC48_DATA_6               (ADC48_DATA_6               ),
    .ADC48_DATA_7               (ADC48_DATA_7               ),
    .ADC48_DATA_8               (ADC48_DATA_8               ),
    .ADC48_DATA_9               (ADC48_DATA_9               ),
    .ADC48_DATA_10              (ADC48_DATA_10              ),
    .ADC48_DATA_11              (ADC48_DATA_11              ),
    .ADC48_DATA_12              (ADC48_DATA_12              ),
    .ADC48_DATA_13              (ADC48_DATA_13              ),
    .ADC48_DATA_14              (ADC48_DATA_14              ),
    .ADC48_DATA_15              (ADC48_DATA_15              ),
    .ADC48_DATA_16              (ADC48_DATA_16              ),
    .ADC48_DATA_17              (ADC48_DATA_17              ),
    .ADC48_DATA_18              (ADC48_DATA_18              ),
    .ADC48_DATA_19              (ADC48_DATA_19              ),
    .ADC48_DATA_20              (ADC48_DATA_20              ),
    .ADC48_DATA_21              (ADC48_DATA_21              ),
    .ADC48_DATA_22              (ADC48_DATA_22              ),
    .ADC48_DATA_23              (ADC48_DATA_23              ),
    .ADC48_DATA_24              (ADC48_DATA_24              ),
    .ADC48_DATA_25              (ADC48_DATA_25              ),
    .ADC48_DATA_26              (ADC48_DATA_26              ),
    .ADC48_DATA_27              (ADC48_DATA_27              ),
    .ADC48_DATA_28              (ADC48_DATA_28              ),
    .ADC48_DATA_29              (ADC48_DATA_29              ),
    .ADC48_DATA_30              (ADC48_DATA_30              ),
    .ADC48_DATA_31              (ADC48_DATA_31              ),
    .ADC48_DATA_32              (ADC48_DATA_32              ),
    .ADC48_DATA_33              (ADC48_DATA_33              ),
    .ADC48_DATA_34              (ADC48_DATA_34              ),
    .ADC48_DATA_35              (ADC48_DATA_35              ),
    .ADC48_DATA_36              (ADC48_DATA_36              ),
    .ADC48_DATA_37              (ADC48_DATA_37              ),
    .ADC48_DATA_38              (ADC48_DATA_38              ),
    .ADC48_DATA_39              (ADC48_DATA_39              ),
    .ADC48_DATA_40              (ADC48_DATA_40              ),
    .ADC48_DATA_41              (ADC48_DATA_41              ),
    .ADC48_DATA_42              (ADC48_DATA_42              ),
    .ADC48_DATA_43              (ADC48_DATA_43              ),
    .ADC48_DATA_44              (ADC48_DATA_44              ),
    .ADC48_DATA_45              (ADC48_DATA_45              ),
    .ADC48_DATA_46              (ADC48_DATA_46              ),
    .ADC48_DATA_47              (ADC48_DATA_47              ),

    .ANA_CLK200M                (ANA_CLK200M                ),
    .ANA_ADC_CLK500M            (ANA_ADC_CLK500M            ),
    .ANA_ADC48_CLK500M          (ANA_ADC48_CLK500M          ),

    .ANA_ADC_DATA_0             (ANA_ADC_DATA_0             ),
    .ANA_ADC_DATA_1             (ANA_ADC_DATA_1             ),
    .ANA_ADC_DATA_2             (ANA_ADC_DATA_2             ),
    .ANA_ADC_DATA_3             (ANA_ADC_DATA_3             ),
    .ANA_ADC_DATA_4             (ANA_ADC_DATA_4             ),
    .ANA_ADC_DATA_5             (ANA_ADC_DATA_5             ),
    .ANA_ADC_DATA_6             (ANA_ADC_DATA_6             ),
    .ANA_ADC_DATA_7             (ANA_ADC_DATA_7             ),
    .ANA_ADC_DATA_8             (ANA_ADC_DATA_8             ),
    .ANA_ADC_DATA_9             (ANA_ADC_DATA_9             ),
    .ANA_ADC_DATA_10            (ANA_ADC_DATA_10            ),
    .ANA_ADC_DATA_11            (ANA_ADC_DATA_11            ),
    .ANA_ADC_DATA_12            (ANA_ADC_DATA_12            ),
    .ANA_ADC_DATA_13            (ANA_ADC_DATA_13            ),
    .ANA_ADC_DATA_14            (ANA_ADC_DATA_14            ),
    .ANA_ADC_DATA_15            (ANA_ADC_DATA_15            ),
    .ANA_ADC_DATA_16            (ANA_ADC_DATA_16            ),
    .ANA_ADC_DATA_17            (ANA_ADC_DATA_17            ),
    .ANA_ADC_DATA_18            (ANA_ADC_DATA_18            ),
    .ANA_ADC_DATA_19            (ANA_ADC_DATA_19            ),
    .ANA_ADC_DATA_20            (ANA_ADC_DATA_20            ),
    .ANA_ADC_DATA_21            (ANA_ADC_DATA_21            ),
    .ANA_ADC_DATA_22            (ANA_ADC_DATA_22            ),
    .ANA_ADC_DATA_23            (ANA_ADC_DATA_23            ),

    .ANA_ADC48_DATA_0           (ANA_ADC48_DATA_0           ),
    .ANA_ADC48_DATA_1           (ANA_ADC48_DATA_1           ),
    .ANA_ADC48_DATA_2           (ANA_ADC48_DATA_2           ),
    .ANA_ADC48_DATA_3           (ANA_ADC48_DATA_3           ),
    .ANA_ADC48_DATA_4           (ANA_ADC48_DATA_4           ),
    .ANA_ADC48_DATA_5           (ANA_ADC48_DATA_5           ),
    .ANA_ADC48_DATA_6           (ANA_ADC48_DATA_6           ),
    .ANA_ADC48_DATA_7           (ANA_ADC48_DATA_7           ),
    .ANA_ADC48_DATA_8           (ANA_ADC48_DATA_8           ),
    .ANA_ADC48_DATA_9           (ANA_ADC48_DATA_9           ),
    .ANA_ADC48_DATA_10          (ANA_ADC48_DATA_10          ),
    .ANA_ADC48_DATA_11          (ANA_ADC48_DATA_11          )
    );

    // crg instantiation
    crg
    u_crg
    (
    .dft_rstnsync_scan_rstn_ctrl(1'b0                       ),
    .dft_rstnsync_scan_rstn     (1'b0                       ),
    .dft_rtl_icg_en             (1'b0                       ),
    .dft_stuck_at_mode          (1'b0                       ),
    .dft_tpi_clk                (1'b0                       ),
    .dft_clkdiv_rstn_ctrl       (1'b0                       ),
    .dft_clkdiv_scan_rstn       (1'b0                       ),
    .dft_scan_en                (1'b0                       ),
    .dft_test_clk_en            (1'b0                       ),
    .ANA_CLK200M                (ANA_CLK200M                ),
    .ANA_ADC_CLK500M            (ANA_ADC_CLK500M            ),
    .ANA_ADC48_CLK500M          (ANA_ADC48_CLK500M          ),
    .rf_96path_en               (rf_96path_en               ),
    .rf_pktctrl_clk_en          (rf_pktctrl_clk_en          ),
    .rf_pktctrl_sw_rstn         (rf_pktctrl_sw_rstn         ),
    .pktctrl_clk                (pktctrl_clk                ),
    .pktctrl_rstn               (pktctrl_rstn               ),
    .clk_200m                   (clk_200m                   ),
    .rstn_200m                  (rstn_200m                  ),
    .adc96_rstn                 (adc96_rstn                 ),
    .adc48_rstn                 (adc48_rstn                 ),
    .RSTN                       (RSTN                       )
    );

    // iopad instantiation
    iopad_top
    u_iopad_top
    (
    .ADC_DATA                   (ADC_DATA                   ),
    .ADC_DATA_VALID             (ADC_DATA_VALID             ),
    .CLK_RD                     (CLK_RD                     ),
    .MDIO_I                     (mdio_out                   ),
    .mdio_oen                   (mdio_oen                   ),
    .RSTN                       (RSTN                       ),
    .MDC                        (MDC                        ),
    .MDIO                       (MDIO                       ),
    .PAD1_ADC_DATA_1            (PAD1_ADC_DATA_1            ),
    .PAD2_ADC_DATA_2            (PAD2_ADC_DATA_2            ),
    .PAD3_ADC_DATA_3            (PAD3_ADC_DATA_3            ),
    .PAD4_ADC_DATA_4            (PAD4_ADC_DATA_4            ),
    .PAD5_ADC_DATA_5            (PAD5_ADC_DATA_5            ),
    .PAD6_ADC_DATA_6            (PAD6_ADC_DATA_6            ),
    .PAD7_ADC_DATA_7            (PAD7_ADC_DATA_7            ),
    .PAD8_ADC_DATA_8            (PAD8_ADC_DATA_8            ),
    .PAD9_ADC_DATA_9            (PAD9_ADC_DATA_9            ),
    .PAD10_ADC_DATA_10          (PAD10_ADC_DATA_10          ),
    .PAD11_ADC_DATA_11          (PAD11_ADC_DATA_11          ),
    .PAD12_ADC_DATA_12          (PAD12_ADC_DATA_12          ),
    .PAD13_ADC_DATA_13          (PAD13_ADC_DATA_13          ),
    .PAD14_ADC_DATA_14          (PAD14_ADC_DATA_14          ),
    .PAD15_ADC_DATA_15          (PAD15_ADC_DATA_15          ),
    .PAD16_ADC_DATA_16          (PAD16_ADC_DATA_16          ),
    .PAD17_ADC_DATA_17          (PAD17_ADC_DATA_17          ),
    .PAD18_ADC_DATA_18          (PAD18_ADC_DATA_18          ),
    .PAD19_ADC_DATA_VALID       (PAD19_ADC_DATA_VALID       ),
    .PAD20_RSTN                 (PAD20_RSTN                 ),
    .PAD21_CLK_RD               (PAD21_CLK_RD               ),
    .PAD22_MDC                  (PAD22_MDC                  ),
    .PAD23_MDIO                 (PAD23_MDIO                 )
    );

    // pktctrl_top instantiation
    pktctrl_top
    u_pktctrl_top
    (
    .pktctrl_clk                (pktctrl_clk                ),
    .pktctrl_rstn               (pktctrl_rstn               ),
    .rf_self_test_mode          (rf_self_test_mode          ),
    .rf_capture_mode            (rf_capture_mode            ),
    .rf_capture_start           (rf_capture_start           ),
    .rf_capture_again           (rf_capture_again           ),
    .rf_96path_en               (rf_96path_en               ),
    .rf_pkt_data_length         (rf_pkt_data_length         ),
    .rf_pkt_idle_length         (rf_pkt_idle_length         ),
    .rf_pktctrl_gap             (rf_pktctrl_gap             ),
    .rf_pktctrl_phase           (rf_pktctrl_phase           ),
    .rf_mdio_data_sel           (rf_mdio_data_sel           ),
    .rf_mdio_memory_addr        (rf_mdio_memory_addr        ),
    .rf_mdio_pkt_data           (rf_mdio_pkt_data           ),
    .ANA_ADC_DATA_0             (ANA_ADC_DATA_0             ),
    .ANA_ADC_DATA_1             (ANA_ADC_DATA_1             ),
    .ANA_ADC_DATA_2             (ANA_ADC_DATA_2             ),
    .ANA_ADC_DATA_3             (ANA_ADC_DATA_3             ),
    .ANA_ADC_DATA_4             (ANA_ADC_DATA_4             ),
    .ANA_ADC_DATA_5             (ANA_ADC_DATA_5             ),
    .ANA_ADC_DATA_6             (ANA_ADC_DATA_6             ),
    .ANA_ADC_DATA_7             (ANA_ADC_DATA_7             ),
    .ANA_ADC_DATA_8             (ANA_ADC_DATA_8             ),
    .ANA_ADC_DATA_9             (ANA_ADC_DATA_9             ),
    .ANA_ADC_DATA_10            (ANA_ADC_DATA_10            ),
    .ANA_ADC_DATA_11            (ANA_ADC_DATA_11            ),
    .ANA_ADC_DATA_12            (ANA_ADC_DATA_12            ),
    .ANA_ADC_DATA_13            (ANA_ADC_DATA_13            ),
    .ANA_ADC_DATA_14            (ANA_ADC_DATA_14            ),
    .ANA_ADC_DATA_15            (ANA_ADC_DATA_15            ),
    .ANA_ADC_DATA_16            (ANA_ADC_DATA_16            ),
    .ANA_ADC_DATA_17            (ANA_ADC_DATA_17            ),
    .ANA_ADC_DATA_18            (ANA_ADC_DATA_18            ),
    .ANA_ADC_DATA_19            (ANA_ADC_DATA_19            ),
    .ANA_ADC_DATA_20            (ANA_ADC_DATA_20            ),
    .ANA_ADC_DATA_21            (ANA_ADC_DATA_21            ),
    .ANA_ADC_DATA_22            (ANA_ADC_DATA_22            ),
    .ANA_ADC_DATA_23            (ANA_ADC_DATA_23            ),
    .ANA_ADC48_DATA_0           (ANA_ADC48_DATA_0           ),
    .ANA_ADC48_DATA_1           (ANA_ADC48_DATA_1           ),
    .ANA_ADC48_DATA_2           (ANA_ADC48_DATA_2           ),
    .ANA_ADC48_DATA_3           (ANA_ADC48_DATA_3           ),
    .ANA_ADC48_DATA_4           (ANA_ADC48_DATA_4           ),
    .ANA_ADC48_DATA_5           (ANA_ADC48_DATA_5           ),
    .ANA_ADC48_DATA_6           (ANA_ADC48_DATA_6           ),
    .ANA_ADC48_DATA_7           (ANA_ADC48_DATA_7           ),
    .ANA_ADC48_DATA_8           (ANA_ADC48_DATA_8           ),
    .ANA_ADC48_DATA_9           (ANA_ADC48_DATA_9           ),
    .ANA_ADC48_DATA_10          (ANA_ADC48_DATA_10          ),
    .ANA_ADC48_DATA_11          (ANA_ADC48_DATA_11          ),
    .CLK_RD                     (CLK_RD                     ),
    .ADC_DATA                   (ADC_DATA                   ),
    .ADC_DATA_VALID             (ADC_DATA_VALID             ),

    //dbg
    .write_info                 (write_info                 ),
    .write_done                 (write_done                 ),
                                                            
    .pkt_ctrl_info              (pkt_ctrl_info              ), 
    .fast_info                  (fast_info                  ), 
    .fast_rd_done               (fast_rd_done               ), 
                                                            
    .fast_main_fsm              (fast_main_fsm              ), 
    .fast_pkt_fsm               (fast_pkt_fsm               ), 
    .idle_cnt                   (idle_cnt                   ), 
    .RD_info                    (RD_info                    )
    );

    // ctrl_sys instantiation
    ctrl_sys
    u_ctrl_sys
    (
    .clk_200m                   (clk_200m                   ),
    .rstn_200m                  (rstn_200m                  ),
    .pktctrl_clk                (pktctrl_clk                ),
    .pktctrl_rstn               (pktctrl_rstn               ),
    .mdio_in                    (MDIO                       ),
    .mdc                        (MDC                        ),
    .mdio_out                   (mdio_out                   ),
    .mdio_oen                   (mdio_oen                   ),
    
    // Digital config register
    .rf_self_test_mode_sync     (rf_self_test_mode          ),
    .rf_capture_mode_sync       (rf_capture_mode            ),
    .rf_capture_start_sync      (rf_capture_start           ),
    .rf_capture_again_sync      (rf_capture_again           ),
    .rf_96path_en_sync          (rf_96path_en               ),
    .rf_pkt_data_length_sync    (rf_pkt_data_length         ),
    .rf_pkt_idle_length_sync    (rf_pkt_idle_length         ),
    .rf_pktctrl_gap_sync        (rf_pktctrl_gap             ),
    .rf_pktctrl_phase_sync      (rf_pktctrl_phase           ),
    .rf_mdio_data_sel_sync      (rf_mdio_data_sel           ),
    .rf_mdio_memory_addr_sync   (rf_mdio_memory_addr        ),
    .rf_mdio_pkt_data           (rf_mdio_pkt_data           ),

    .rf_pktctrl_clk_en          (rf_pktctrl_clk_en          ),
    .rf_pktctrl_sw_rstn         (rf_pktctrl_sw_rstn         ),

    .capture_enable             (capture_enable             ),
    .capture_start              (capture_start              ),

    .capture_mode               (capture_mode               ),
    .capture_max_addr           (capture_max_addr           ),
    .pre_trigger_num            (pre_trigger_num            ),

    .trigger_pattern0           (trigger_pattern0           ),
    .trigger_pattern1           (trigger_pattern1           ),
    .trigger_mode0              (trigger_mode0              ),
    .trigger_mode1              (trigger_mode1              ),
    .trigger_mode2              (trigger_mode2              ),
    .trigger_mode3              (trigger_mode3              ),
    .trigger_mode4              (trigger_mode4              ),
    .trigger_mode5              (trigger_mode5              ),
    .trigger_logic0             (trigger_logic0             ),
    .trigger_logic1             (trigger_logic1             ),
    .store_mode                 (store_mode                 ),

    .read_start_addr            (read_start_addr            ),
    .tri_addr                   (tri_addr                   ),
    .capture_done_rd            (capture_done_rd            ),
    .capture_done               (capture_done               ),

    .tri_succeed_cnt_overflow_mode(tri_succeed_cnt_overflow_mode),
    .tri_succeed_cnt_clr        (tri_succeed_cnt_clr        ),
    .tri_succeed_cnt            (tri_succeed_cnt            ),

    .capture_rd_en              (capture_rd_en              ),
    .capture_rd_addr            (capture_rd_addr            ),
    .capture_rd_data0           (capture_rd_data0           ),
    .capture_rd_data1           (capture_rd_data1           )
    );

    dbg_top
    u_dbg_top
    (
    .wr_clk                     (pktctrl_clk                ),
    .wr_rst_n                   (pktctrl_rstn               ),
    .rd_clk                     (clk_200m                   ),
    .rd_rst_n                   (rstn_200m                  ),
                                                            
    .write_info                 (write_info                 ), 
    .write_done                 (write_done                 ), 
                                                            
    .pkt_ctrl_info              (pkt_ctrl_info              ), 
    .fast_info                  (fast_info                  ), 
    .fast_rd_done               (fast_rd_done               ), 
                                                            
    .fast_main_fsm              (fast_main_fsm              ), 
    .fast_pkt_fsm               (fast_pkt_fsm               ), 
    .idle_cnt                   (idle_cnt                   ), 
    .RD_info                    (RD_info                    ), 
                                                            
    .tri_succeed                (tri_succeed                ), //TODO TODO
    .tri_data                   (tri_data                   ),
    .tri_data_vld               (tri_data_vld               ),
                                                            
    .capture_enable             (capture_enable             ),
    .capture_start              (capture_start              ),

    .capture_mode               (capture_mode               ),
    .capture_max_addr           (capture_max_addr           ),
    .pre_trigger_num            (pre_trigger_num            ),

    .trigger_pattern0           (trigger_pattern0           ),
    .trigger_pattern1           (trigger_pattern1           ),
    .trigger_mode0              (trigger_mode0              ),
    .trigger_mode1              (trigger_mode1              ),
    .trigger_mode2              (trigger_mode2              ),
    .trigger_mode3              (trigger_mode3              ),
    .trigger_mode4              (trigger_mode4              ),
    .trigger_mode5              (trigger_mode5              ),
    .trigger_logic0             (trigger_logic0             ),
    .trigger_logic1             (trigger_logic1             ),
    .store_mode                 (store_mode                 ),

    .read_start_addr            (read_start_addr            ),
    .tri_addr                   (tri_addr                   ),
    .capture_done_rd            (capture_done_rd            ),
    .capture_done               (capture_done               ),

    .tri_succeed_cnt_overflow_mode(tri_succeed_cnt_overflow_mode),
    .tri_succeed_cnt_clr        (tri_succeed_cnt_clr        ),
    .tri_succeed_cnt            (tri_succeed_cnt            ),

    .capture_rd_en              (capture_rd_en              ),
    .capture_rd_addr            (capture_rd_addr            ),
    .capture_rd_data0           (capture_rd_data0           ),
    .capture_rd_data1           (capture_rd_data1           )
    );

endmodule
