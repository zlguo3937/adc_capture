module design_C ( input_tc , net_c1_a1, net_b1_c1, net_c1_a2, net_c1_a3, net_b3_c1_a2,
                  output_tc, net_b2_c2, net_c2_a2, net_b1_c2, net_c2_a3, net_a3_b1_c2,
                  inout_tc , net_b1_c3, net_b2_c3, net_c3_a1_b2
                );
    input   input_tc ,
            net_c1_a1, net_b1_c1,
            net_c1_a2, net_c1_a3, net_b3_c1_a2;
    output  output_tc,
            net_b2_c2, net_c2_a2,
            net_b1_c2, net_c2_a3, net_a3_b1_c2;
    inout   inout_tc , net_b1_c3,
            net_b2_c3, net_c3_a1_b2;

    //assign ...
    //always ...

endmodule

