module ANALOG_WRAPPER
(
    output  wire    CLK200M,
    output  wire    CLK500M
);

endmodule
