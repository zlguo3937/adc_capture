# Created by MC2 : Version 2012.02.00.d on 2024/05/10, 15:14:14

#*********************************************************************************************************************/
# Software       : TSMC MEMORY COMPILER tsn28hpcpd127spsram_2012.02.00.d.180a						*/
# Technology     : TSMC 28nm CMOS LOGIC High Performance Compact Mobile Computing Plus 1P10M HKMG CU_ELK 0.9V				*/
#  Memory Type    : TSMC 28nm High Performance Compact Mobile Computing Plus Single Port SRAM with d127 bit cell HVT periphery */
# Library Name   : ts1n28hpcphvtb16384x36m8sso (user specify : TS1N28HPCPHVTB16384X36M8SSO)				*/
# Library Version: 180a												*/
# Generated Time : 2024/05/10, 15:14:06										*/
#*********************************************************************************************************************/
#															*/
# STATEMENT OF USE													*/
#															*/
# This information contains confidential and proprietary information of TSMC.					*/
# No part of this information may be reproduced, transmitted, transcribed,						*/
# stored in a retrieval system, or translated into any human or computer						*/
# language, in any form or by any means, electronic, mechanical, magnetic,						*/
# optical, chemical, manual, or otherwise, without the prior written permission					*/
# of TSMC. This information was prepared for informational purpose and is for					*/
# use by TSMC's customers only. TSMC reserves the right to make changes in the					*/
# information at any time and without notice.									*/
#															*/
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS1N28HPCPHVTB16384X36M8SSO
	CLASS BLOCK ;
	FOREIGN TS1N28HPCPHVTB16384X36M8SSO 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 653.535 BY 186.370 ;
	SYMMETRY X Y ;
	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 95.670 653.535 95.820 ;
			LAYER M3 ;
			RECT 653.355 95.670 653.535 95.820 ;
			LAYER M1 ;
			RECT 653.355 95.670 653.535 95.820 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[0]

	PIN A[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 85.420 653.535 85.570 ;
			LAYER M3 ;
			RECT 653.355 85.420 653.535 85.570 ;
			LAYER M2 ;
			RECT 653.355 85.420 653.535 85.570 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[10]

	PIN A[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 98.110 653.535 98.260 ;
			LAYER M1 ;
			RECT 653.355 98.110 653.535 98.260 ;
			LAYER M2 ;
			RECT 653.355 98.110 653.535 98.260 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[11]

	PIN A[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 97.720 653.535 97.870 ;
			LAYER M1 ;
			RECT 653.355 97.720 653.535 97.870 ;
			LAYER M3 ;
			RECT 653.355 97.720 653.535 97.870 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[12]

	PIN A[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 96.060 653.535 96.210 ;
			LAYER M2 ;
			RECT 653.355 96.060 653.535 96.210 ;
			LAYER M3 ;
			RECT 653.355 96.060 653.535 96.210 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[13]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 94.010 653.535 94.160 ;
			LAYER M3 ;
			RECT 653.355 94.010 653.535 94.160 ;
			LAYER M1 ;
			RECT 653.355 94.010 653.535 94.160 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 93.620 653.535 93.770 ;
			LAYER M3 ;
			RECT 653.355 93.620 653.535 93.770 ;
			LAYER M2 ;
			RECT 653.355 93.620 653.535 93.770 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 89.520 653.535 89.670 ;
			LAYER M2 ;
			RECT 653.355 89.520 653.535 89.670 ;
			LAYER M3 ;
			RECT 653.355 89.520 653.535 89.670 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 87.860 653.535 88.010 ;
			LAYER M3 ;
			RECT 653.355 87.860 653.535 88.010 ;
			LAYER M1 ;
			RECT 653.355 87.860 653.535 88.010 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 87.470 653.535 87.620 ;
			LAYER M2 ;
			RECT 653.355 87.470 653.535 87.620 ;
			LAYER M1 ;
			RECT 653.355 87.470 653.535 87.620 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 91.960 653.535 92.110 ;
			LAYER M2 ;
			RECT 653.355 91.960 653.535 92.110 ;
			LAYER M1 ;
			RECT 653.355 91.960 653.535 92.110 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 91.570 653.535 91.720 ;
			LAYER M3 ;
			RECT 653.355 91.570 653.535 91.720 ;
			LAYER M1 ;
			RECT 653.355 91.570 653.535 91.720 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 89.910 653.535 90.060 ;
			LAYER M1 ;
			RECT 653.355 89.910 653.535 90.060 ;
			LAYER M3 ;
			RECT 653.355 89.910 653.535 90.060 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 85.810 653.535 85.960 ;
			LAYER M1 ;
			RECT 653.355 85.810 653.535 85.960 ;
			LAYER M3 ;
			RECT 653.355 85.810 653.535 85.960 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[9]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 99.770 653.535 99.920 ;
			LAYER M3 ;
			RECT 653.355 99.770 653.535 99.920 ;
			LAYER M2 ;
			RECT 653.355 99.770 653.535 99.920 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.115300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.228300 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.515900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.249900 LAYER M2 ;
		ANTENNAMAXAREACAR 10.191100 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.732500 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 11.091100 LAYER M3 ;
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 100.400 653.535 100.550 ;
			LAYER M2 ;
			RECT 653.355 100.400 653.535 100.550 ;
			LAYER M3 ;
			RECT 653.355 100.400 653.535 100.550 ;
		END
		ANTENNAGATEAREA 2.013900 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 3.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 5.372500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.331500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA1 ;
		ANTENNAGATEAREA 2.013900 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 2.694600 LAYER M2 ;
		ANTENNAMAXAREACAR 33.912400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.292500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.097200 LAYER VIA2 ;
		ANTENNAGATEAREA 2.013900 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 2.754400 LAYER M3 ;
		ANTENNAMAXAREACAR 35.107800 LAYER M3 ;
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 4.315 653.535 4.465 ;
			LAYER M1 ;
			RECT 653.355 4.315 653.535 4.465 ;
			LAYER M2 ;
			RECT 653.355 4.315 653.535 4.465 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[0]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 50.715 653.535 50.865 ;
			LAYER M2 ;
			RECT 653.355 50.715 653.535 50.865 ;
			LAYER M3 ;
			RECT 653.355 50.715 653.535 50.865 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 55.355 653.535 55.505 ;
			LAYER M2 ;
			RECT 653.355 55.355 653.535 55.505 ;
			LAYER M3 ;
			RECT 653.355 55.355 653.535 55.505 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 59.995 653.535 60.145 ;
			LAYER M2 ;
			RECT 653.355 59.995 653.535 60.145 ;
			LAYER M3 ;
			RECT 653.355 59.995 653.535 60.145 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 64.635 653.535 64.785 ;
			LAYER M2 ;
			RECT 653.355 64.635 653.535 64.785 ;
			LAYER M1 ;
			RECT 653.355 64.635 653.535 64.785 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 69.275 653.535 69.425 ;
			LAYER M2 ;
			RECT 653.355 69.275 653.535 69.425 ;
			LAYER M3 ;
			RECT 653.355 69.275 653.535 69.425 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 73.915 653.535 74.065 ;
			LAYER M2 ;
			RECT 653.355 73.915 653.535 74.065 ;
			LAYER M1 ;
			RECT 653.355 73.915 653.535 74.065 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 76.235 653.535 76.385 ;
			LAYER M1 ;
			RECT 653.355 76.235 653.535 76.385 ;
			LAYER M3 ;
			RECT 653.355 76.235 653.535 76.385 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 78.555 653.535 78.705 ;
			LAYER M3 ;
			RECT 653.355 78.555 653.535 78.705 ;
			LAYER M1 ;
			RECT 653.355 78.555 653.535 78.705 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 107.275 653.535 107.425 ;
			LAYER M2 ;
			RECT 653.355 107.275 653.535 107.425 ;
			LAYER M1 ;
			RECT 653.355 107.275 653.535 107.425 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 109.595 653.535 109.745 ;
			LAYER M2 ;
			RECT 653.355 109.595 653.535 109.745 ;
			LAYER M3 ;
			RECT 653.355 109.595 653.535 109.745 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[19]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 8.955 653.535 9.105 ;
			LAYER M1 ;
			RECT 653.355 8.955 653.535 9.105 ;
			LAYER M3 ;
			RECT 653.355 8.955 653.535 9.105 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[1]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 114.235 653.535 114.385 ;
			LAYER M1 ;
			RECT 653.355 114.235 653.535 114.385 ;
			LAYER M3 ;
			RECT 653.355 114.235 653.535 114.385 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 118.875 653.535 119.025 ;
			LAYER M2 ;
			RECT 653.355 118.875 653.535 119.025 ;
			LAYER M3 ;
			RECT 653.355 118.875 653.535 119.025 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 123.515 653.535 123.665 ;
			LAYER M2 ;
			RECT 653.355 123.515 653.535 123.665 ;
			LAYER M1 ;
			RECT 653.355 123.515 653.535 123.665 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 128.155 653.535 128.305 ;
			LAYER M3 ;
			RECT 653.355 128.155 653.535 128.305 ;
			LAYER M2 ;
			RECT 653.355 128.155 653.535 128.305 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 132.795 653.535 132.945 ;
			LAYER M3 ;
			RECT 653.355 132.795 653.535 132.945 ;
			LAYER M2 ;
			RECT 653.355 132.795 653.535 132.945 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 137.435 653.535 137.585 ;
			LAYER M3 ;
			RECT 653.355 137.435 653.535 137.585 ;
			LAYER M1 ;
			RECT 653.355 137.435 653.535 137.585 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 142.075 653.535 142.225 ;
			LAYER M1 ;
			RECT 653.355 142.075 653.535 142.225 ;
			LAYER M3 ;
			RECT 653.355 142.075 653.535 142.225 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 146.715 653.535 146.865 ;
			LAYER M1 ;
			RECT 653.355 146.715 653.535 146.865 ;
			LAYER M2 ;
			RECT 653.355 146.715 653.535 146.865 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 151.355 653.535 151.505 ;
			LAYER M3 ;
			RECT 653.355 151.355 653.535 151.505 ;
			LAYER M2 ;
			RECT 653.355 151.355 653.535 151.505 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 155.995 653.535 156.145 ;
			LAYER M1 ;
			RECT 653.355 155.995 653.535 156.145 ;
			LAYER M2 ;
			RECT 653.355 155.995 653.535 156.145 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[29]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 13.595 653.535 13.745 ;
			LAYER M3 ;
			RECT 653.355 13.595 653.535 13.745 ;
			LAYER M1 ;
			RECT 653.355 13.595 653.535 13.745 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[2]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 160.635 653.535 160.785 ;
			LAYER M3 ;
			RECT 653.355 160.635 653.535 160.785 ;
			LAYER M2 ;
			RECT 653.355 160.635 653.535 160.785 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 165.275 653.535 165.425 ;
			LAYER M3 ;
			RECT 653.355 165.275 653.535 165.425 ;
			LAYER M1 ;
			RECT 653.355 165.275 653.535 165.425 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[31]

	PIN D[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 169.915 653.535 170.065 ;
			LAYER M1 ;
			RECT 653.355 169.915 653.535 170.065 ;
			LAYER M2 ;
			RECT 653.355 169.915 653.535 170.065 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[32]

	PIN D[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 174.555 653.535 174.705 ;
			LAYER M3 ;
			RECT 653.355 174.555 653.535 174.705 ;
			LAYER M1 ;
			RECT 653.355 174.555 653.535 174.705 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[33]

	PIN D[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 179.195 653.535 179.345 ;
			LAYER M1 ;
			RECT 653.355 179.195 653.535 179.345 ;
			LAYER M2 ;
			RECT 653.355 179.195 653.535 179.345 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[34]

	PIN D[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 183.835 653.535 183.985 ;
			LAYER M2 ;
			RECT 653.355 183.835 653.535 183.985 ;
			LAYER M1 ;
			RECT 653.355 183.835 653.535 183.985 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[35]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 18.235 653.535 18.385 ;
			LAYER M3 ;
			RECT 653.355 18.235 653.535 18.385 ;
			LAYER M1 ;
			RECT 653.355 18.235 653.535 18.385 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 22.875 653.535 23.025 ;
			LAYER M2 ;
			RECT 653.355 22.875 653.535 23.025 ;
			LAYER M3 ;
			RECT 653.355 22.875 653.535 23.025 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 27.515 653.535 27.665 ;
			LAYER M3 ;
			RECT 653.355 27.515 653.535 27.665 ;
			LAYER M1 ;
			RECT 653.355 27.515 653.535 27.665 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 32.155 653.535 32.305 ;
			LAYER M2 ;
			RECT 653.355 32.155 653.535 32.305 ;
			LAYER M1 ;
			RECT 653.355 32.155 653.535 32.305 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 36.795 653.535 36.945 ;
			LAYER M2 ;
			RECT 653.355 36.795 653.535 36.945 ;
			LAYER M3 ;
			RECT 653.355 36.795 653.535 36.945 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 41.435 653.535 41.585 ;
			LAYER M2 ;
			RECT 653.355 41.435 653.535 41.585 ;
			LAYER M1 ;
			RECT 653.355 41.435 653.535 41.585 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 46.075 653.535 46.225 ;
			LAYER M2 ;
			RECT 653.355 46.075 653.535 46.225 ;
			LAYER M1 ;
			RECT 653.355 46.075 653.535 46.225 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[9]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 5.325 653.535 5.475 ;
			LAYER M2 ;
			RECT 653.355 5.325 653.535 5.475 ;
			LAYER M1 ;
			RECT 653.355 5.325 653.535 5.475 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[0]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 51.725 653.535 51.875 ;
			LAYER M1 ;
			RECT 653.355 51.725 653.535 51.875 ;
			LAYER M3 ;
			RECT 653.355 51.725 653.535 51.875 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 56.365 653.535 56.515 ;
			LAYER M2 ;
			RECT 653.355 56.365 653.535 56.515 ;
			LAYER M3 ;
			RECT 653.355 56.365 653.535 56.515 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 61.005 653.535 61.155 ;
			LAYER M3 ;
			RECT 653.355 61.005 653.535 61.155 ;
			LAYER M2 ;
			RECT 653.355 61.005 653.535 61.155 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 65.645 653.535 65.795 ;
			LAYER M2 ;
			RECT 653.355 65.645 653.535 65.795 ;
			LAYER M3 ;
			RECT 653.355 65.645 653.535 65.795 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 70.285 653.535 70.435 ;
			LAYER M3 ;
			RECT 653.355 70.285 653.535 70.435 ;
			LAYER M1 ;
			RECT 653.355 70.285 653.535 70.435 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 74.925 653.535 75.075 ;
			LAYER M1 ;
			RECT 653.355 74.925 653.535 75.075 ;
			LAYER M3 ;
			RECT 653.355 74.925 653.535 75.075 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 77.245 653.535 77.395 ;
			LAYER M1 ;
			RECT 653.355 77.245 653.535 77.395 ;
			LAYER M3 ;
			RECT 653.355 77.245 653.535 77.395 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 79.565 653.535 79.715 ;
			LAYER M2 ;
			RECT 653.355 79.565 653.535 79.715 ;
			LAYER M1 ;
			RECT 653.355 79.565 653.535 79.715 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 108.285 653.535 108.435 ;
			LAYER M2 ;
			RECT 653.355 108.285 653.535 108.435 ;
			LAYER M1 ;
			RECT 653.355 108.285 653.535 108.435 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 110.605 653.535 110.755 ;
			LAYER M2 ;
			RECT 653.355 110.605 653.535 110.755 ;
			LAYER M3 ;
			RECT 653.355 110.605 653.535 110.755 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[19]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 9.965 653.535 10.115 ;
			LAYER M2 ;
			RECT 653.355 9.965 653.535 10.115 ;
			LAYER M1 ;
			RECT 653.355 9.965 653.535 10.115 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[1]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 115.245 653.535 115.395 ;
			LAYER M3 ;
			RECT 653.355 115.245 653.535 115.395 ;
			LAYER M2 ;
			RECT 653.355 115.245 653.535 115.395 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 119.885 653.535 120.035 ;
			LAYER M3 ;
			RECT 653.355 119.885 653.535 120.035 ;
			LAYER M2 ;
			RECT 653.355 119.885 653.535 120.035 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 124.525 653.535 124.675 ;
			LAYER M1 ;
			RECT 653.355 124.525 653.535 124.675 ;
			LAYER M2 ;
			RECT 653.355 124.525 653.535 124.675 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 129.165 653.535 129.315 ;
			LAYER M3 ;
			RECT 653.355 129.165 653.535 129.315 ;
			LAYER M2 ;
			RECT 653.355 129.165 653.535 129.315 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 133.805 653.535 133.955 ;
			LAYER M1 ;
			RECT 653.355 133.805 653.535 133.955 ;
			LAYER M3 ;
			RECT 653.355 133.805 653.535 133.955 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 138.445 653.535 138.595 ;
			LAYER M1 ;
			RECT 653.355 138.445 653.535 138.595 ;
			LAYER M3 ;
			RECT 653.355 138.445 653.535 138.595 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 143.085 653.535 143.235 ;
			LAYER M1 ;
			RECT 653.355 143.085 653.535 143.235 ;
			LAYER M3 ;
			RECT 653.355 143.085 653.535 143.235 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 147.725 653.535 147.875 ;
			LAYER M2 ;
			RECT 653.355 147.725 653.535 147.875 ;
			LAYER M1 ;
			RECT 653.355 147.725 653.535 147.875 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 152.365 653.535 152.515 ;
			LAYER M2 ;
			RECT 653.355 152.365 653.535 152.515 ;
			LAYER M1 ;
			RECT 653.355 152.365 653.535 152.515 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 157.005 653.535 157.155 ;
			LAYER M1 ;
			RECT 653.355 157.005 653.535 157.155 ;
			LAYER M3 ;
			RECT 653.355 157.005 653.535 157.155 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[29]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 14.605 653.535 14.755 ;
			LAYER M3 ;
			RECT 653.355 14.605 653.535 14.755 ;
			LAYER M1 ;
			RECT 653.355 14.605 653.535 14.755 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[2]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 161.645 653.535 161.795 ;
			LAYER M1 ;
			RECT 653.355 161.645 653.535 161.795 ;
			LAYER M2 ;
			RECT 653.355 161.645 653.535 161.795 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 166.285 653.535 166.435 ;
			LAYER M1 ;
			RECT 653.355 166.285 653.535 166.435 ;
			LAYER M3 ;
			RECT 653.355 166.285 653.535 166.435 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[31]

	PIN Q[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 170.925 653.535 171.075 ;
			LAYER M1 ;
			RECT 653.355 170.925 653.535 171.075 ;
			LAYER M3 ;
			RECT 653.355 170.925 653.535 171.075 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[32]

	PIN Q[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 175.565 653.535 175.715 ;
			LAYER M3 ;
			RECT 653.355 175.565 653.535 175.715 ;
			LAYER M2 ;
			RECT 653.355 175.565 653.535 175.715 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[33]

	PIN Q[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 180.205 653.535 180.355 ;
			LAYER M2 ;
			RECT 653.355 180.205 653.535 180.355 ;
			LAYER M3 ;
			RECT 653.355 180.205 653.535 180.355 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[34]

	PIN Q[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 184.845 653.535 184.995 ;
			LAYER M2 ;
			RECT 653.355 184.845 653.535 184.995 ;
			LAYER M3 ;
			RECT 653.355 184.845 653.535 184.995 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[35]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 19.245 653.535 19.395 ;
			LAYER M1 ;
			RECT 653.355 19.245 653.535 19.395 ;
			LAYER M3 ;
			RECT 653.355 19.245 653.535 19.395 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 23.885 653.535 24.035 ;
			LAYER M2 ;
			RECT 653.355 23.885 653.535 24.035 ;
			LAYER M3 ;
			RECT 653.355 23.885 653.535 24.035 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 28.525 653.535 28.675 ;
			LAYER M1 ;
			RECT 653.355 28.525 653.535 28.675 ;
			LAYER M3 ;
			RECT 653.355 28.525 653.535 28.675 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 33.165 653.535 33.315 ;
			LAYER M1 ;
			RECT 653.355 33.165 653.535 33.315 ;
			LAYER M3 ;
			RECT 653.355 33.165 653.535 33.315 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 37.805 653.535 37.955 ;
			LAYER M1 ;
			RECT 653.355 37.805 653.535 37.955 ;
			LAYER M2 ;
			RECT 653.355 37.805 653.535 37.955 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 42.445 653.535 42.595 ;
			LAYER M1 ;
			RECT 653.355 42.445 653.535 42.595 ;
			LAYER M2 ;
			RECT 653.355 42.445 653.535 42.595 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 653.355 47.085 653.535 47.235 ;
			LAYER M2 ;
			RECT 653.355 47.085 653.535 47.235 ;
			LAYER M1 ;
			RECT 653.355 47.085 653.535 47.235 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[9]

	PIN SD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 81.145 653.535 81.295 ;
			LAYER M1 ;
			RECT 653.355 81.145 653.535 81.295 ;
			LAYER M3 ;
			RECT 653.355 81.145 653.535 81.295 ;
		END
		ANTENNAGATEAREA 0.051000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.839700 LAYER M1 ;
		ANTENNAMAXAREACAR 9.087800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.585600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.051000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.499900 LAYER M2 ;
		ANTENNAMAXAREACAR 48.990700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.878400 LAYER VIA2 ;
		ANTENNAGATEAREA 0.051000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.590600 LAYER M3 ;
		ANTENNAMAXAREACAR 48.990700 LAYER M3 ;
	END SD

	PIN SLP
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 653.355 81.860 653.535 82.010 ;
			LAYER M1 ;
			RECT 653.355 81.860 653.535 82.010 ;
			LAYER M3 ;
			RECT 653.355 81.860 653.535 82.010 ;
		END
		ANTENNAGATEAREA 0.027000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.172400 LAYER M1 ;
		ANTENNAMAXAREACAR 8.260000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.433300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.027000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.269000 LAYER M2 ;
		ANTENNAMAXAREACAR 48.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.027000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.564300 LAYER M3 ;
		ANTENNAMAXAREACAR 48.814800 LAYER M3 ;
	END SLP

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.000 2.555 653.145 2.885 ;
			LAYER M4 ;
			RECT 0.000 7.195 653.145 7.525 ;
			LAYER M4 ;
			RECT 0.000 11.835 653.145 12.165 ;
			LAYER M4 ;
			RECT 0.000 16.475 653.145 16.805 ;
			LAYER M4 ;
			RECT 0.000 21.115 653.145 21.445 ;
			LAYER M4 ;
			RECT 0.000 25.755 653.145 26.085 ;
			LAYER M4 ;
			RECT 0.000 30.395 653.145 30.725 ;
			LAYER M4 ;
			RECT 0.000 35.035 653.145 35.365 ;
			LAYER M4 ;
			RECT 0.000 39.675 653.145 40.005 ;
			LAYER M4 ;
			RECT 0.000 44.315 653.145 44.645 ;
			LAYER M4 ;
			RECT 0.000 48.955 653.145 49.285 ;
			LAYER M4 ;
			RECT 0.000 53.595 653.145 53.925 ;
			LAYER M4 ;
			RECT 0.000 58.235 653.145 58.565 ;
			LAYER M4 ;
			RECT 0.000 62.875 653.145 63.205 ;
			LAYER M4 ;
			RECT 0.000 67.515 653.145 67.845 ;
			LAYER M4 ;
			RECT 0.000 72.155 653.145 72.485 ;
			LAYER M4 ;
			RECT 0.000 76.795 653.535 77.125 ;
			LAYER M4 ;
			RECT 0.000 81.435 653.535 81.765 ;
			LAYER M4 ;
			RECT 0.000 91.755 653.535 92.325 ;
			LAYER M4 ;
			RECT 0.000 92.455 653.535 93.025 ;
			LAYER M4 ;
			RECT 0.000 99.435 653.535 100.005 ;
			LAYER M4 ;
			RECT 0.000 103.195 653.535 103.525 ;
			LAYER M4 ;
			RECT 0.000 107.835 653.535 108.165 ;
			LAYER M4 ;
			RECT 0.000 112.475 653.145 112.805 ;
			LAYER M4 ;
			RECT 0.000 117.115 653.145 117.445 ;
			LAYER M4 ;
			RECT 0.000 121.755 653.145 122.085 ;
			LAYER M4 ;
			RECT 0.000 126.395 653.145 126.725 ;
			LAYER M4 ;
			RECT 0.000 131.035 653.145 131.365 ;
			LAYER M4 ;
			RECT 0.000 135.675 653.145 136.005 ;
			LAYER M4 ;
			RECT 0.000 140.315 653.145 140.645 ;
			LAYER M4 ;
			RECT 0.000 144.955 653.145 145.285 ;
			LAYER M4 ;
			RECT 0.000 149.595 653.145 149.925 ;
			LAYER M4 ;
			RECT 0.000 154.235 653.145 154.565 ;
			LAYER M4 ;
			RECT 0.000 158.875 653.145 159.205 ;
			LAYER M4 ;
			RECT 0.000 163.515 653.145 163.845 ;
			LAYER M4 ;
			RECT 0.000 168.155 653.145 168.485 ;
			LAYER M4 ;
			RECT 0.000 172.795 653.145 173.125 ;
			LAYER M4 ;
			RECT 0.000 177.435 653.145 177.765 ;
			LAYER M4 ;
			RECT 0.000 182.075 653.145 182.405 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.000 3.965 653.145 4.345 ;
			LAYER M4 ;
			RECT 0.000 8.605 653.145 8.985 ;
			LAYER M4 ;
			RECT 0.000 13.245 653.145 13.625 ;
			LAYER M4 ;
			RECT 0.000 17.885 653.145 18.265 ;
			LAYER M4 ;
			RECT 0.000 22.525 653.145 22.905 ;
			LAYER M4 ;
			RECT 0.000 27.165 653.145 27.545 ;
			LAYER M4 ;
			RECT 0.000 31.805 653.145 32.185 ;
			LAYER M4 ;
			RECT 0.000 36.445 653.145 36.825 ;
			LAYER M4 ;
			RECT 0.000 41.085 653.145 41.465 ;
			LAYER M4 ;
			RECT 0.000 45.725 653.145 46.105 ;
			LAYER M4 ;
			RECT 0.000 50.365 653.145 50.745 ;
			LAYER M4 ;
			RECT 0.000 55.005 653.145 55.385 ;
			LAYER M4 ;
			RECT 0.000 59.645 653.145 60.025 ;
			LAYER M4 ;
			RECT 0.000 64.285 653.145 64.665 ;
			LAYER M4 ;
			RECT 0.000 68.925 653.145 69.305 ;
			LAYER M4 ;
			RECT 0.000 73.565 653.145 73.945 ;
			LAYER M4 ;
			RECT 0.000 78.205 653.535 78.585 ;
			LAYER M4 ;
			RECT 0.000 82.845 653.535 83.225 ;
			LAYER M4 ;
			RECT 0.000 90.355 653.535 90.925 ;
			LAYER M4 ;
			RECT 0.000 91.055 653.535 91.625 ;
			LAYER M4 ;
			RECT 0.000 93.385 653.535 93.955 ;
			LAYER M4 ;
			RECT 0.000 104.605 653.535 104.985 ;
			LAYER M4 ;
			RECT 0.000 109.245 653.535 109.625 ;
			LAYER M4 ;
			RECT 0.000 113.885 653.145 114.265 ;
			LAYER M4 ;
			RECT 0.000 118.525 653.145 118.905 ;
			LAYER M4 ;
			RECT 0.000 123.165 653.145 123.545 ;
			LAYER M4 ;
			RECT 0.000 127.805 653.145 128.185 ;
			LAYER M4 ;
			RECT 0.000 132.445 653.145 132.825 ;
			LAYER M4 ;
			RECT 0.000 137.085 653.145 137.465 ;
			LAYER M4 ;
			RECT 0.000 141.725 653.145 142.105 ;
			LAYER M4 ;
			RECT 0.000 146.365 653.145 146.745 ;
			LAYER M4 ;
			RECT 0.000 151.005 653.145 151.385 ;
			LAYER M4 ;
			RECT 0.000 155.645 653.145 156.025 ;
			LAYER M4 ;
			RECT 0.000 160.285 653.145 160.665 ;
			LAYER M4 ;
			RECT 0.000 164.925 653.145 165.305 ;
			LAYER M4 ;
			RECT 0.000 169.565 653.145 169.945 ;
			LAYER M4 ;
			RECT 0.000 174.205 653.145 174.585 ;
			LAYER M4 ;
			RECT 0.000 178.845 653.145 179.225 ;
			LAYER M4 ;
			RECT 0.000 183.485 653.145 183.865 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 653.355 83.370 653.535 83.520 ;
			LAYER M3 ;
			RECT 653.355 83.370 653.535 83.520 ;
			LAYER M2 ;
			RECT 653.355 83.370 653.535 83.520 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.445400 LAYER M2 ;
		ANTENNAMAXAREACAR 16.888300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 17.788300 LAYER M3 ;
	END WEB

	OBS
		# Promoted blockages
		LAYER M1 ;
		RECT 653.355 185.055 653.535 186.370 ;
		LAYER M3 ;
		RECT 653.355 185.075 653.535 186.370 ;
		LAYER VIA3 ;
		RECT 653.355 185.075 653.535 186.370 ;
		LAYER M1 ;
		RECT 653.355 143.295 653.535 146.655 ;
		LAYER M1 ;
		RECT 653.355 61.215 653.535 64.575 ;
		LAYER M3 ;
		RECT 653.355 60.225 653.535 60.925 ;
		LAYER VIA3 ;
		RECT 653.355 60.225 653.535 60.925 ;
		LAYER M2 ;
		RECT 653.355 60.225 653.535 60.925 ;
		LAYER M1 ;
		RECT 653.355 27.725 653.535 28.465 ;
		LAYER M2 ;
		RECT 653.355 33.395 653.535 36.715 ;
		LAYER M3 ;
		RECT 653.355 33.395 653.535 36.715 ;
		LAYER M2 ;
		RECT 653.355 37.025 653.535 37.725 ;
		LAYER M3 ;
		RECT 653.355 27.745 653.535 28.445 ;
		LAYER VIA3 ;
		RECT 653.355 27.745 653.535 28.445 ;
		LAYER M2 ;
		RECT 653.355 24.115 653.535 27.435 ;
		LAYER M3 ;
		RECT 653.355 24.115 653.535 27.435 ;
		LAYER VIA3 ;
		RECT 653.355 24.115 653.535 27.435 ;
		LAYER M3 ;
		RECT 653.355 61.235 653.535 64.555 ;
		LAYER M2 ;
		RECT 653.355 64.865 653.535 65.565 ;
		LAYER M1 ;
		RECT 653.355 65.855 653.535 69.215 ;
		LAYER M1 ;
		RECT 653.355 24.095 653.535 27.455 ;
		LAYER M1 ;
		RECT 653.355 56.575 653.535 59.935 ;
		LAYER M1 ;
		RECT 653.355 60.205 653.535 60.945 ;
		LAYER M3 ;
		RECT 653.355 64.865 653.535 65.565 ;
		LAYER M3 ;
		RECT 653.355 78.785 653.535 79.485 ;
		LAYER M1 ;
		RECT 653.355 92.170 653.535 93.560 ;
		LAYER M2 ;
		RECT 653.355 91.800 653.535 91.880 ;
		LAYER M1 ;
		RECT 653.355 142.285 653.535 143.025 ;
		LAYER M1 ;
		RECT 653.355 120.095 653.535 123.455 ;
		LAYER M3 ;
		RECT 653.355 120.115 653.535 123.435 ;
		LAYER M3 ;
		RECT 653.355 142.305 653.535 143.005 ;
		LAYER M2 ;
		RECT 653.355 142.305 653.535 143.005 ;
		LAYER M2 ;
		RECT 653.355 128.385 653.535 129.085 ;
		LAYER M3 ;
		RECT 653.355 128.385 653.535 129.085 ;
		LAYER M1 ;
		RECT 653.355 123.725 653.535 124.465 ;
		LAYER VIA3 ;
		RECT 653.355 128.385 653.535 129.085 ;
		LAYER M3 ;
		RECT 653.355 56.595 653.535 59.915 ;
		LAYER VIA3 ;
		RECT 653.355 56.595 653.535 59.915 ;
		LAYER VIA3 ;
		RECT 653.355 50.945 653.535 51.645 ;
		LAYER M3 ;
		RECT 653.355 51.955 653.535 55.275 ;
		LAYER VIA3 ;
		RECT 653.355 51.955 653.535 55.275 ;
		LAYER M1 ;
		RECT 653.355 50.925 653.535 51.665 ;
		LAYER M3 ;
		RECT 653.355 46.305 653.535 47.005 ;
		LAYER M2 ;
		RECT 653.355 46.305 653.535 47.005 ;
		LAYER VIA3 ;
		RECT 653.355 46.305 653.535 47.005 ;
		LAYER M1 ;
		RECT 653.355 46.285 653.535 47.025 ;
		LAYER M2 ;
		RECT 653.355 47.315 653.535 50.635 ;
		LAYER M3 ;
		RECT 653.355 42.675 653.535 45.995 ;
		LAYER VIA3 ;
		RECT 653.355 42.675 653.535 45.995 ;
		LAYER M2 ;
		RECT 653.355 42.675 653.535 45.995 ;
		LAYER M1 ;
		RECT 653.355 42.655 653.535 46.015 ;
		LAYER M1 ;
		RECT 653.355 55.565 653.535 56.305 ;
		LAYER M3 ;
		RECT 653.355 55.585 653.535 56.285 ;
		LAYER VIA3 ;
		RECT 653.355 55.585 653.535 56.285 ;
		LAYER M2 ;
		RECT 653.355 55.585 653.535 56.285 ;
		LAYER M3 ;
		RECT 653.355 47.315 653.535 50.635 ;
		LAYER VIA3 ;
		RECT 653.355 47.315 653.535 50.635 ;
		LAYER M1 ;
		RECT 653.355 47.295 653.535 50.655 ;
		LAYER M2 ;
		RECT 653.355 28.755 653.535 32.075 ;
		LAYER M1 ;
		RECT 653.355 32.365 653.535 33.105 ;
		LAYER VIA3 ;
		RECT 653.355 33.395 653.535 36.715 ;
		LAYER M3 ;
		RECT 653.355 28.755 653.535 32.075 ;
		LAYER VIA3 ;
		RECT 653.355 28.755 653.535 32.075 ;
		LAYER M1 ;
		RECT 653.355 33.375 653.535 36.735 ;
		LAYER M1 ;
		RECT 653.355 37.005 653.535 37.745 ;
		LAYER M3 ;
		RECT 653.355 37.025 653.535 37.725 ;
		LAYER VIA3 ;
		RECT 653.355 37.025 653.535 37.725 ;
		LAYER M1 ;
		RECT 653.355 38.015 653.535 41.375 ;
		LAYER M1 ;
		RECT 653.355 28.735 653.535 32.095 ;
		LAYER M2 ;
		RECT 653.355 32.385 653.535 33.085 ;
		LAYER M3 ;
		RECT 653.355 32.385 653.535 33.085 ;
		LAYER VIA3 ;
		RECT 653.355 32.385 653.535 33.085 ;
		LAYER M2 ;
		RECT 653.355 185.075 653.535 186.370 ;
		LAYER M1 ;
		RECT 653.355 180.415 653.535 183.775 ;
		LAYER VIA3 ;
		RECT 653.355 180.435 653.535 183.755 ;
		LAYER M1 ;
		RECT 653.355 184.045 653.535 184.785 ;
		LAYER M2 ;
		RECT 653.355 184.065 653.535 184.765 ;
		LAYER M2 ;
		RECT 653.355 180.435 653.535 183.755 ;
		LAYER M3 ;
		RECT 653.355 180.435 653.535 183.755 ;
		LAYER M3 ;
		RECT 653.355 184.065 653.535 184.765 ;
		LAYER VIA3 ;
		RECT 653.355 184.065 653.535 184.765 ;
		LAYER M2 ;
		RECT 653.355 152.595 653.535 155.915 ;
		LAYER M1 ;
		RECT 653.355 152.575 653.535 155.935 ;
		LAYER VIA3 ;
		RECT 653.355 156.225 653.535 156.925 ;
		LAYER M2 ;
		RECT 653.355 156.225 653.535 156.925 ;
		LAYER M2 ;
		RECT 653.355 165.505 653.535 166.205 ;
		LAYER M3 ;
		RECT 653.355 170.145 653.535 170.845 ;
		LAYER VIA3 ;
		RECT 653.355 170.145 653.535 170.845 ;
		LAYER VIA3 ;
		RECT 653.355 165.505 653.535 166.205 ;
		LAYER M3 ;
		RECT 653.355 165.505 653.535 166.205 ;
		LAYER M2 ;
		RECT 653.355 171.155 653.535 174.475 ;
		LAYER M3 ;
		RECT 653.355 171.155 653.535 174.475 ;
		LAYER M1 ;
		RECT 653.355 170.125 653.535 170.865 ;
		LAYER M2 ;
		RECT 653.355 174.785 653.535 175.485 ;
		LAYER VIA3 ;
		RECT 653.355 174.785 653.535 175.485 ;
		LAYER M1 ;
		RECT 653.355 171.135 653.535 174.495 ;
		LAYER M3 ;
		RECT 653.355 174.785 653.535 175.485 ;
		LAYER VIA3 ;
		RECT 653.355 171.155 653.535 174.475 ;
		LAYER M2 ;
		RECT 653.355 160.865 653.535 161.565 ;
		LAYER M3 ;
		RECT 653.355 160.865 653.535 161.565 ;
		LAYER M2 ;
		RECT 653.355 157.235 653.535 160.555 ;
		LAYER M3 ;
		RECT 653.355 157.235 653.535 160.555 ;
		LAYER VIA3 ;
		RECT 653.355 160.865 653.535 161.565 ;
		LAYER VIA3 ;
		RECT 653.355 157.235 653.535 160.555 ;
		LAYER M3 ;
		RECT 653.355 161.875 653.535 165.195 ;
		LAYER VIA3 ;
		RECT 653.355 161.875 653.535 165.195 ;
		LAYER M2 ;
		RECT 653.355 161.875 653.535 165.195 ;
		LAYER M1 ;
		RECT 653.355 161.855 653.535 165.215 ;
		LAYER M2 ;
		RECT 653.355 166.515 653.535 169.835 ;
		LAYER M3 ;
		RECT 653.355 166.515 653.535 169.835 ;
		LAYER VIA3 ;
		RECT 653.355 166.515 653.535 169.835 ;
		LAYER M2 ;
		RECT 653.355 170.145 653.535 170.845 ;
		LAYER VIA3 ;
		RECT 653.355 75.155 653.535 76.155 ;
		LAYER M2 ;
		RECT 653.355 75.155 653.535 76.155 ;
		LAYER M3 ;
		RECT 653.355 75.155 653.535 76.155 ;
		LAYER M3 ;
		RECT 653.355 74.145 653.535 74.845 ;
		LAYER VIA3 ;
		RECT 653.355 74.145 653.535 74.845 ;
		LAYER M3 ;
		RECT 653.355 79.795 653.535 81.065 ;
		LAYER VIA3 ;
		RECT 653.355 79.795 653.535 81.065 ;
		LAYER M2 ;
		RECT 653.355 81.375 653.535 81.780 ;
		LAYER M2 ;
		RECT 653.355 70.515 653.535 73.835 ;
		LAYER M1 ;
		RECT 653.355 82.070 653.535 83.310 ;
		LAYER M3 ;
		RECT 653.355 81.375 653.535 81.780 ;
		LAYER M2 ;
		RECT 653.355 86.040 653.535 87.390 ;
		LAYER M1 ;
		RECT 653.355 86.020 653.535 87.410 ;
		LAYER M2 ;
		RECT 653.355 85.650 653.535 85.730 ;
		LAYER M1 ;
		RECT 653.355 85.630 653.535 85.750 ;
		LAYER VIA3 ;
		RECT 653.355 85.650 653.535 85.730 ;
		LAYER M3 ;
		RECT 653.355 175.795 653.535 179.115 ;
		LAYER M1 ;
		RECT 653.355 160.845 653.535 161.585 ;
		LAYER M1 ;
		RECT 653.355 174.765 653.535 175.505 ;
		LAYER M3 ;
		RECT 653.355 179.425 653.535 180.125 ;
		LAYER VIA3 ;
		RECT 653.355 179.425 653.535 180.125 ;
		LAYER M1 ;
		RECT 653.355 175.775 653.535 179.135 ;
		LAYER M2 ;
		RECT 653.355 179.425 653.535 180.125 ;
		LAYER M1 ;
		RECT 653.355 179.405 653.535 180.145 ;
		LAYER M2 ;
		RECT 653.355 175.795 653.535 179.115 ;
		LAYER VIA3 ;
		RECT 653.355 175.795 653.535 179.115 ;
		LAYER M3 ;
		RECT 653.355 152.595 653.535 155.915 ;
		LAYER VIA3 ;
		RECT 653.355 152.595 653.535 155.915 ;
		LAYER M3 ;
		RECT 653.355 156.225 653.535 156.925 ;
		LAYER M2 ;
		RECT 653.355 65.875 653.535 69.195 ;
		LAYER M1 ;
		RECT 653.355 70.495 653.535 73.855 ;
		LAYER M2 ;
		RECT 653.355 89.750 653.535 89.830 ;
		LAYER M1 ;
		RECT 653.355 89.730 653.535 89.850 ;
		LAYER M3 ;
		RECT 653.355 151.585 653.535 152.285 ;
		LAYER VIA3 ;
		RECT 653.355 151.585 653.535 152.285 ;
		LAYER M3 ;
		RECT 653.355 147.955 653.535 151.275 ;
		LAYER VIA3 ;
		RECT 653.355 147.955 653.535 151.275 ;
		LAYER M1 ;
		RECT 653.355 151.565 653.535 152.305 ;
		LAYER M2 ;
		RECT 653.355 151.585 653.535 152.285 ;
		LAYER M1 ;
		RECT 653.355 134.015 653.535 137.375 ;
		LAYER M1 ;
		RECT 653.355 133.005 653.535 133.745 ;
		LAYER M2 ;
		RECT 653.355 97.950 653.535 98.030 ;
		LAYER M3 ;
		RECT 653.355 146.945 653.535 147.645 ;
		LAYER M3 ;
		RECT 653.355 143.315 653.535 146.635 ;
		LAYER M2 ;
		RECT 653.355 143.315 653.535 146.635 ;
		LAYER VIA3 ;
		RECT 653.355 143.315 653.535 146.635 ;
		LAYER M2 ;
		RECT 653.355 146.945 653.535 147.645 ;
		LAYER VIA3 ;
		RECT 653.355 146.945 653.535 147.645 ;
		LAYER M1 ;
		RECT 653.355 147.935 653.535 151.295 ;
		LAYER M1 ;
		RECT 653.355 146.925 653.535 147.665 ;
		LAYER M1 ;
		RECT 653.355 138.655 653.535 142.015 ;
		LAYER M2 ;
		RECT 653.355 147.955 653.535 151.275 ;
		LAYER VIA3 ;
		RECT 653.355 142.305 653.535 143.005 ;
		LAYER M3 ;
		RECT 653.355 138.675 653.535 141.995 ;
		LAYER M3 ;
		RECT 653.355 134.035 653.535 137.355 ;
		LAYER VIA3 ;
		RECT 653.355 134.035 653.535 137.355 ;
		LAYER VIA3 ;
		RECT 653.355 137.665 653.535 138.365 ;
		LAYER M3 ;
		RECT 653.355 137.665 653.535 138.365 ;
		LAYER VIA3 ;
		RECT 653.355 133.025 653.535 133.725 ;
		LAYER M2 ;
		RECT 653.355 137.665 653.535 138.365 ;
		LAYER M1 ;
		RECT 653.355 137.645 653.535 138.385 ;
		LAYER M2 ;
		RECT 653.355 134.035 653.535 137.355 ;
		LAYER M2 ;
		RECT 653.355 133.025 653.535 133.725 ;
		LAYER M3 ;
		RECT 653.355 133.025 653.535 133.725 ;
		LAYER M2 ;
		RECT 653.355 138.675 653.535 141.995 ;
		LAYER M2 ;
		RECT 653.355 129.395 653.535 132.715 ;
		LAYER VIA3 ;
		RECT 653.355 123.745 653.535 124.445 ;
		LAYER M3 ;
		RECT 653.355 115.475 653.535 118.795 ;
		LAYER M2 ;
		RECT 653.355 98.340 653.535 99.690 ;
		LAYER M3 ;
		RECT 653.355 100.000 653.535 100.320 ;
		LAYER VIA3 ;
		RECT 653.355 100.000 653.535 100.320 ;
		LAYER M2 ;
		RECT 653.355 100.000 653.535 100.320 ;
		LAYER VIA3 ;
		RECT 653.355 98.340 653.535 99.690 ;
		LAYER M1 ;
		RECT 653.355 108.495 653.535 109.535 ;
		LAYER M2 ;
		RECT 653.355 107.505 653.535 108.205 ;
		LAYER M3 ;
		RECT 653.355 107.505 653.535 108.205 ;
		LAYER M1 ;
		RECT 653.355 107.485 653.535 108.225 ;
		LAYER M1 ;
		RECT 653.355 100.610 653.535 107.215 ;
		LAYER M3 ;
		RECT 653.355 98.340 653.535 99.690 ;
		LAYER VIA3 ;
		RECT 653.355 93.850 653.535 93.930 ;
		LAYER M1 ;
		RECT 653.355 99.980 653.535 100.340 ;
		LAYER VIA3 ;
		RECT 653.355 138.675 653.535 141.995 ;
		LAYER M3 ;
		RECT 653.355 129.395 653.535 132.715 ;
		LAYER VIA3 ;
		RECT 653.355 129.395 653.535 132.715 ;
		LAYER M1 ;
		RECT 653.355 129.375 653.535 132.735 ;
		LAYER M1 ;
		RECT 653.355 128.365 653.535 129.105 ;
		LAYER M2 ;
		RECT 653.355 100.630 653.535 107.195 ;
		LAYER VIA3 ;
		RECT 653.355 107.505 653.535 108.205 ;
		LAYER M1 ;
		RECT 653.355 115.455 653.535 118.815 ;
		LAYER VIA3 ;
		RECT 653.355 119.105 653.535 119.805 ;
		LAYER M3 ;
		RECT 653.355 100.630 653.535 107.195 ;
		LAYER VIA3 ;
		RECT 653.355 100.630 653.535 107.195 ;
		LAYER M1 ;
		RECT 653.355 119.085 653.535 119.825 ;
		LAYER M1 ;
		RECT 653.355 74.125 653.535 74.865 ;
		LAYER M2 ;
		RECT 653.355 74.145 653.535 74.845 ;
		LAYER M1 ;
		RECT 653.355 75.135 653.535 76.175 ;
		LAYER M1 ;
		RECT 653.355 124.735 653.535 128.095 ;
		LAYER M2 ;
		RECT 653.355 124.755 653.535 128.075 ;
		LAYER M3 ;
		RECT 653.355 124.755 653.535 128.075 ;
		LAYER M2 ;
		RECT 653.355 123.745 653.535 124.445 ;
		LAYER VIA3 ;
		RECT 653.355 124.755 653.535 128.075 ;
		LAYER M3 ;
		RECT 653.355 123.745 653.535 124.445 ;
		LAYER M2 ;
		RECT 653.355 119.105 653.535 119.805 ;
		LAYER M3 ;
		RECT 653.355 119.105 653.535 119.805 ;
		LAYER M2 ;
		RECT 653.355 120.115 653.535 123.435 ;
		LAYER VIA3 ;
		RECT 653.355 120.115 653.535 123.435 ;
		LAYER M2 ;
		RECT 653.355 76.465 653.535 77.165 ;
		LAYER M3 ;
		RECT 653.355 76.465 653.535 77.165 ;
		LAYER M2 ;
		RECT 653.355 77.475 653.535 78.475 ;
		LAYER M3 ;
		RECT 653.355 77.475 653.535 78.475 ;
		LAYER M1 ;
		RECT 653.355 78.765 653.535 79.505 ;
		LAYER VIA3 ;
		RECT 653.355 78.785 653.535 79.485 ;
		LAYER M2 ;
		RECT 653.355 78.785 653.535 79.485 ;
		LAYER M1 ;
		RECT 653.355 93.830 653.535 93.950 ;
		LAYER M2 ;
		RECT 653.355 93.850 653.535 93.930 ;
		LAYER M3 ;
		RECT 653.355 93.850 653.535 93.930 ;
		LAYER VIA3 ;
		RECT 653.355 92.190 653.535 93.540 ;
		LAYER M1 ;
		RECT 653.355 97.930 653.535 98.050 ;
		LAYER M3 ;
		RECT 653.355 91.800 653.535 91.880 ;
		LAYER M1 ;
		RECT 653.355 77.455 653.535 78.495 ;
		LAYER M1 ;
		RECT 653.355 98.320 653.535 99.710 ;
		LAYER M2 ;
		RECT 653.355 110.835 653.535 114.155 ;
		LAYER VIA3 ;
		RECT 653.355 110.835 653.535 114.155 ;
		LAYER M2 ;
		RECT 653.355 79.795 653.535 81.065 ;
		LAYER M1 ;
		RECT 653.355 79.775 653.535 81.085 ;
		LAYER M2 ;
		RECT 653.355 90.140 653.535 91.490 ;
		LAYER M1 ;
		RECT 653.355 90.120 653.535 91.510 ;
		LAYER M3 ;
		RECT 653.355 90.140 653.535 91.490 ;
		LAYER VIA3 ;
		RECT 653.355 90.140 653.535 91.490 ;
		LAYER M2 ;
		RECT 653.355 94.240 653.535 95.590 ;
		LAYER M3 ;
		RECT 653.355 94.240 653.535 95.590 ;
		LAYER VIA3 ;
		RECT 653.355 91.800 653.535 91.880 ;
		LAYER M2 ;
		RECT 653.355 51.955 653.535 55.275 ;
		LAYER M1 ;
		RECT 653.355 51.935 653.535 55.295 ;
		LAYER M3 ;
		RECT 653.355 50.945 653.535 51.645 ;
		LAYER M2 ;
		RECT 653.355 50.945 653.535 51.645 ;
		LAYER M3 ;
		RECT 653.355 38.035 653.535 41.355 ;
		LAYER M2 ;
		RECT 653.355 38.035 653.535 41.355 ;
		LAYER VIA3 ;
		RECT 653.355 38.035 653.535 41.355 ;
		LAYER M2 ;
		RECT 653.355 41.665 653.535 42.365 ;
		LAYER VIA3 ;
		RECT 653.355 41.665 653.535 42.365 ;
		LAYER M3 ;
		RECT 653.355 41.665 653.535 42.365 ;
		LAYER M1 ;
		RECT 653.355 41.645 653.535 42.385 ;
		LAYER M3 ;
		RECT 653.355 65.875 653.535 69.195 ;
		LAYER VIA3 ;
		RECT 653.355 65.875 653.535 69.195 ;
		LAYER M3 ;
		RECT 653.355 70.515 653.535 73.835 ;
		LAYER VIA3 ;
		RECT 653.355 70.515 653.535 73.835 ;
		LAYER M3 ;
		RECT 653.355 97.950 653.535 98.030 ;
		LAYER M2 ;
		RECT 653.355 95.900 653.535 95.980 ;
		LAYER VIA3 ;
		RECT 653.355 94.240 653.535 95.590 ;
		LAYER M1 ;
		RECT 653.355 95.880 653.535 96.000 ;
		LAYER M1 ;
		RECT 653.355 94.220 653.535 95.610 ;
		LAYER VIA3 ;
		RECT 653.355 97.950 653.535 98.030 ;
		LAYER M3 ;
		RECT 653.355 88.090 653.535 89.440 ;
		LAYER M1 ;
		RECT 653.355 76.445 653.535 77.185 ;
		LAYER VIA3 ;
		RECT 653.355 76.465 653.535 77.165 ;
		LAYER M2 ;
		RECT 653.355 69.505 653.535 70.205 ;
		LAYER M3 ;
		RECT 653.355 69.505 653.535 70.205 ;
		LAYER VIA3 ;
		RECT 653.355 69.505 653.535 70.205 ;
		LAYER M1 ;
		RECT 653.355 69.485 653.535 70.225 ;
		LAYER M2 ;
		RECT 653.355 82.090 653.535 83.290 ;
		LAYER M3 ;
		RECT 653.355 82.090 653.535 83.290 ;
		LAYER VIA3 ;
		RECT 653.355 82.090 653.535 83.290 ;
		LAYER VIA3 ;
		RECT 653.355 77.475 653.535 78.475 ;
		LAYER VIA3 ;
		RECT 653.355 81.375 653.535 81.780 ;
		LAYER M1 ;
		RECT 653.355 81.355 653.535 81.800 ;
		LAYER M1 ;
		RECT 653.355 88.070 653.535 89.460 ;
		LAYER M3 ;
		RECT 653.355 89.750 653.535 89.830 ;
		LAYER VIA3 ;
		RECT 653.355 89.750 653.535 89.830 ;
		LAYER M1 ;
		RECT 653.355 91.780 653.535 91.900 ;
		LAYER M3 ;
		RECT 653.355 92.190 653.535 93.540 ;
		LAYER M2 ;
		RECT 653.355 92.190 653.535 93.540 ;
		LAYER M2 ;
		RECT 653.355 88.090 653.535 89.440 ;
		LAYER VIA3 ;
		RECT 653.355 88.090 653.535 89.440 ;
		LAYER VIA3 ;
		RECT 653.355 86.040 653.535 87.390 ;
		LAYER M1 ;
		RECT 653.355 87.680 653.535 87.800 ;
		LAYER M2 ;
		RECT 653.355 83.600 653.535 85.340 ;
		LAYER VIA3 ;
		RECT 653.355 83.600 653.535 85.340 ;
		LAYER M1 ;
		RECT 653.355 83.580 653.535 85.360 ;
		LAYER M3 ;
		RECT 653.355 83.600 653.535 85.340 ;
		LAYER M3 ;
		RECT 653.355 85.650 653.535 85.730 ;
		LAYER M2 ;
		RECT 653.355 96.290 653.535 97.640 ;
		LAYER M3 ;
		RECT 653.355 96.290 653.535 97.640 ;
		LAYER VIA3 ;
		RECT 653.355 96.290 653.535 97.640 ;
		LAYER M1 ;
		RECT 653.355 96.270 653.535 97.660 ;
		LAYER M3 ;
		RECT 653.355 95.900 653.535 95.980 ;
		LAYER VIA3 ;
		RECT 653.355 95.900 653.535 95.980 ;
		LAYER M2 ;
		RECT 653.355 87.700 653.535 87.780 ;
		LAYER M3 ;
		RECT 653.355 87.700 653.535 87.780 ;
		LAYER VIA3 ;
		RECT 653.355 87.700 653.535 87.780 ;
		LAYER M3 ;
		RECT 653.355 86.040 653.535 87.390 ;
		LAYER VIA3 ;
		RECT 653.355 115.475 653.535 118.795 ;
		LAYER M3 ;
		RECT 653.355 114.465 653.535 115.165 ;
		LAYER VIA3 ;
		RECT 653.355 114.465 653.535 115.165 ;
		LAYER M1 ;
		RECT 653.355 114.445 653.535 115.185 ;
		LAYER M2 ;
		RECT 653.355 114.465 653.535 115.165 ;
		LAYER M2 ;
		RECT 653.355 115.475 653.535 118.795 ;
		LAYER M1 ;
		RECT 653.355 110.815 653.535 114.175 ;
		LAYER M3 ;
		RECT 653.355 110.835 653.535 114.155 ;
		LAYER M2 ;
		RECT 653.355 109.825 653.535 110.525 ;
		LAYER M3 ;
		RECT 653.355 109.825 653.535 110.525 ;
		LAYER VIA3 ;
		RECT 653.355 109.825 653.535 110.525 ;
		LAYER M1 ;
		RECT 653.355 109.805 653.535 110.545 ;
		LAYER M2 ;
		RECT 653.355 108.515 653.535 109.515 ;
		LAYER M3 ;
		RECT 653.355 108.515 653.535 109.515 ;
		LAYER VIA3 ;
		RECT 653.355 108.515 653.535 109.515 ;
		LAYER M1 ;
		RECT 653.355 166.495 653.535 169.855 ;
		LAYER M1 ;
		RECT 653.355 165.485 653.535 166.225 ;
		LAYER M1 ;
		RECT 653.355 157.215 653.535 160.575 ;
		LAYER M1 ;
		RECT 653.355 156.205 653.535 156.945 ;
		LAYER M1 ;
		RECT 653.355 9.165 653.535 9.905 ;
		LAYER M2 ;
		RECT 653.355 9.185 653.535 9.885 ;
		LAYER M3 ;
		RECT 653.355 9.185 653.535 9.885 ;
		LAYER VIA3 ;
		RECT 653.355 9.185 653.535 9.885 ;
		LAYER M2 ;
		RECT 653.355 5.555 653.535 8.875 ;
		LAYER M3 ;
		RECT 653.355 5.555 653.535 8.875 ;
		LAYER M2 ;
		RECT 653.355 10.195 653.535 13.515 ;
		LAYER M3 ;
		RECT 653.355 10.195 653.535 13.515 ;
		LAYER M1 ;
		RECT 653.355 10.175 653.535 13.535 ;
		LAYER VIA3 ;
		RECT 653.355 5.555 653.535 8.875 ;
		LAYER VIA3 ;
		RECT 653.355 64.865 653.535 65.565 ;
		LAYER M1 ;
		RECT 653.355 13.805 653.535 14.545 ;
		LAYER VIA3 ;
		RECT 653.355 10.195 653.535 13.515 ;
		LAYER M2 ;
		RECT 653.355 18.465 653.535 19.165 ;
		LAYER M2 ;
		RECT 653.355 14.835 653.535 18.155 ;
		LAYER M3 ;
		RECT 653.355 14.835 653.535 18.155 ;
		LAYER M2 ;
		RECT 653.355 13.825 653.535 14.525 ;
		LAYER VIA3 ;
		RECT 653.355 14.835 653.535 18.155 ;
		LAYER M1 ;
		RECT 653.355 14.815 653.535 18.175 ;
		LAYER M3 ;
		RECT 653.355 18.465 653.535 19.165 ;
		LAYER M3 ;
		RECT 653.355 13.825 653.535 14.525 ;
		LAYER VIA3 ;
		RECT 653.355 13.825 653.535 14.525 ;
		LAYER M1 ;
		RECT 653.355 64.845 653.535 65.585 ;
		LAYER M2 ;
		RECT 653.355 23.105 653.535 23.805 ;
		LAYER M1 ;
		RECT 653.355 23.085 653.535 23.825 ;
		LAYER M1 ;
		RECT 653.355 19.455 653.535 22.815 ;
		LAYER M2 ;
		RECT 653.355 27.745 653.535 28.445 ;
		LAYER M1 ;
		RECT 653.355 4.525 653.535 5.265 ;
		LAYER M1 ;
		RECT 653.355 0.000 653.535 4.255 ;
		LAYER M2 ;
		RECT 653.355 0.000 653.535 4.235 ;
		LAYER VIA3 ;
		RECT 653.355 4.545 653.535 5.245 ;
		LAYER M4 ;
		RECT 0.000 78.585 653.535 79.580 ;
		LAYER M4 ;
		RECT 0.000 143.910 653.145 144.955 ;
		LAYER M4 ;
		RECT 0.000 151.385 653.145 152.380 ;
		LAYER M4 ;
		RECT 0.000 157.830 653.145 158.875 ;
		LAYER M4 ;
		RECT 0.000 156.025 653.145 157.020 ;
		LAYER M4 ;
		RECT 0.000 134.630 653.145 135.675 ;
		LAYER M4 ;
		RECT 0.000 67.845 653.145 68.925 ;
		LAYER M3 ;
		RECT 0.000 0.000 653.355 186.370 ;
		LAYER M4 ;
		RECT 0.000 159.205 653.145 160.285 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 653.355 186.370 ;
		LAYER M4 ;
		RECT 0.000 160.665 653.145 161.660 ;
		LAYER M4 ;
		RECT 0.000 179.225 653.145 180.220 ;
		LAYER M4 ;
		RECT 0.000 171.750 653.145 172.795 ;
		LAYER M4 ;
		RECT 0.000 169.945 653.145 170.940 ;
		LAYER M4 ;
		RECT 0.000 142.105 653.145 143.100 ;
		LAYER M4 ;
		RECT 0.000 140.645 653.145 141.725 ;
		LAYER M4 ;
		RECT 0.000 154.565 653.145 155.645 ;
		LAYER M4 ;
		RECT 0.000 149.925 653.145 151.005 ;
		LAYER M4 ;
		RECT 0.000 148.550 653.145 149.595 ;
		LAYER M4 ;
		RECT 0.000 153.190 653.145 154.235 ;
		LAYER M4 ;
		RECT 229.605 100.005 247.735 101.540 ;
		LAYER M4 ;
		RECT 195.045 100.585 229.605 101.540 ;
		LAYER M4 ;
		RECT 0.000 137.465 653.145 138.460 ;
		LAYER M4 ;
		RECT 0.000 100.005 1.315 101.540 ;
		LAYER M4 ;
		RECT 0.000 165.305 653.145 166.300 ;
		LAYER M4 ;
		RECT 0.000 163.845 653.145 164.925 ;
		LAYER M4 ;
		RECT 0.000 177.765 653.145 178.845 ;
		LAYER M4 ;
		RECT 0.000 176.390 653.145 177.435 ;
		LAYER M4 ;
		RECT 0.000 174.585 653.145 175.580 ;
		LAYER M4 ;
		RECT 0.000 173.125 653.145 174.205 ;
		LAYER M4 ;
		RECT 353.515 100.585 373.495 101.540 ;
		LAYER M4 ;
		RECT 318.255 100.585 352.815 101.540 ;
		LAYER M4 ;
		RECT 0.000 111.430 653.145 112.475 ;
		LAYER M4 ;
		RECT 318.255 100.005 373.495 100.585 ;
		LAYER M4 ;
		RECT 317.555 100.005 318.255 101.540 ;
		LAYER M4 ;
		RECT 0.000 146.745 653.145 147.740 ;
		LAYER M4 ;
		RECT 0.000 145.285 653.145 146.365 ;
		LAYER M4 ;
		RECT 89.805 100.585 123.825 101.540 ;
		LAYER M4 ;
		RECT 124.525 100.585 159.085 101.540 ;
		LAYER M4 ;
		RECT 159.785 100.585 194.345 101.540 ;
		LAYER M4 ;
		RECT 89.265 100.005 159.085 100.585 ;
		LAYER M4 ;
		RECT 1.315 100.585 35.875 101.540 ;
		LAYER M4 ;
		RECT 1.315 100.005 71.135 100.585 ;
		LAYER M4 ;
		RECT 0.000 136.005 653.145 137.085 ;
		LAYER M4 ;
		RECT 0.000 139.270 653.145 140.315 ;
		LAYER M3 ;
		RECT 653.355 0.000 653.535 4.235 ;
		LAYER VIA3 ;
		RECT 653.355 0.000 653.535 4.235 ;
		LAYER M2 ;
		RECT 653.355 4.545 653.535 5.245 ;
		LAYER M3 ;
		RECT 653.355 4.545 653.535 5.245 ;
		LAYER M4 ;
		RECT 0.000 162.470 653.145 163.515 ;
		LAYER M4 ;
		RECT 0.000 1.510 653.145 2.555 ;
		LAYER M4 ;
		RECT 0.000 2.885 653.145 3.965 ;
		LAYER M4 ;
		RECT 0.000 4.345 653.145 5.340 ;
		LAYER M4 ;
		RECT 0.000 6.150 653.145 7.195 ;
		LAYER M1 ;
		RECT 653.355 5.535 653.535 8.895 ;
		LAYER VIA3 ;
		RECT 653.355 18.465 653.535 19.165 ;
		LAYER M2 ;
		RECT 653.355 19.475 653.535 22.795 ;
		LAYER M1 ;
		RECT 653.355 18.445 653.535 19.185 ;
		LAYER M3 ;
		RECT 653.355 19.475 653.535 22.795 ;
		LAYER VIA3 ;
		RECT 653.355 19.475 653.535 22.795 ;
		LAYER M3 ;
		RECT 653.355 23.105 653.535 23.805 ;
		LAYER VIA3 ;
		RECT 653.355 23.105 653.535 23.805 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 653.535 186.370 ;
		LAYER M4 ;
		RECT 0.000 168.485 653.145 169.565 ;
		LAYER M4 ;
		RECT 0.000 181.030 653.145 182.075 ;
		LAYER M4 ;
		RECT 0.000 182.405 653.145 183.485 ;
		LAYER M1 ;
		RECT 0.000 0.000 653.355 186.370 ;
		LAYER M4 ;
		RECT 0.000 183.865 653.145 184.860 ;
		LAYER M4 ;
		RECT 0.000 167.110 653.145 168.155 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 653.535 186.370 ;
		LAYER M2 ;
		RECT 0.000 0.000 653.355 186.370 ;
		LAYER M2 ;
		RECT 653.355 61.235 653.535 64.555 ;
		LAYER VIA3 ;
		RECT 653.355 61.235 653.535 64.555 ;
		LAYER M2 ;
		RECT 653.355 56.595 653.535 59.915 ;
		LAYER M4 ;
		RECT 653.145 100.005 653.535 103.195 ;
		LAYER M4 ;
		RECT 635.675 93.025 653.535 93.385 ;
		LAYER M4 ;
		RECT 0.000 93.955 653.535 99.435 ;
		LAYER M4 ;
		RECT 0.000 84.535 653.535 90.355 ;
		LAYER M4 ;
		RECT 71.135 100.005 89.265 101.540 ;
		LAYER M4 ;
		RECT 159.085 100.005 159.785 101.540 ;
		LAYER M4 ;
		RECT 0.000 132.825 653.145 133.820 ;
		LAYER M4 ;
		RECT 0.000 123.545 653.145 124.540 ;
		LAYER M4 ;
		RECT 0.000 102.150 636.335 103.195 ;
		LAYER M4 ;
		RECT 0.000 103.525 653.535 104.605 ;
		LAYER M4 ;
		RECT 0.000 116.070 653.145 117.115 ;
		LAYER M4 ;
		RECT 0.000 117.445 653.145 118.525 ;
		LAYER M4 ;
		RECT 0.000 114.265 653.145 115.260 ;
		LAYER M4 ;
		RECT 0.000 112.805 653.145 113.885 ;
		LAYER M4 ;
		RECT 636.335 104.985 653.535 106.150 ;
		LAYER M4 ;
		RECT 0.000 122.085 653.145 123.165 ;
		LAYER M4 ;
		RECT 0.000 120.710 653.145 121.755 ;
		LAYER M4 ;
		RECT 636.335 101.540 653.145 103.195 ;
		LAYER M4 ;
		RECT 373.495 100.005 653.145 101.540 ;
		LAYER M4 ;
		RECT 247.735 100.005 317.555 100.585 ;
		LAYER M4 ;
		RECT 0.000 131.365 653.145 132.445 ;
		LAYER M4 ;
		RECT 0.000 128.185 653.145 129.180 ;
		LAYER M4 ;
		RECT 0.000 126.725 653.145 127.805 ;
		LAYER M4 ;
		RECT 0.000 125.350 653.145 126.395 ;
		LAYER M4 ;
		RECT 0.000 129.990 653.145 131.035 ;
		LAYER M4 ;
		RECT 0.000 104.985 636.335 105.980 ;
		LAYER M4 ;
		RECT 0.000 106.790 653.535 107.835 ;
		LAYER M4 ;
		RECT 0.000 108.165 653.535 109.245 ;
		LAYER M4 ;
		RECT 0.000 118.905 653.145 119.900 ;
		LAYER M4 ;
		RECT 0.000 109.625 653.535 110.620 ;
		LAYER M4 ;
		RECT 36.575 100.585 71.135 101.540 ;
		LAYER M4 ;
		RECT 248.275 100.585 282.295 101.540 ;
		LAYER M4 ;
		RECT 282.995 100.585 317.555 101.540 ;
		LAYER M4 ;
		RECT 159.785 100.005 229.605 100.585 ;
		LAYER M4 ;
		RECT 0.000 52.550 653.145 53.595 ;
		LAYER M4 ;
		RECT 0.000 53.925 653.145 55.005 ;
		LAYER M4 ;
		RECT 0.000 55.385 653.145 56.380 ;
		LAYER M4 ;
		RECT 0.000 64.665 653.145 65.660 ;
		LAYER M4 ;
		RECT 0.000 63.205 653.145 64.285 ;
		LAYER M4 ;
		RECT 0.000 61.830 653.145 62.875 ;
		LAYER M4 ;
		RECT 0.000 60.025 653.145 61.020 ;
		LAYER M4 ;
		RECT 0.000 58.565 653.145 59.645 ;
		LAYER M4 ;
		RECT 0.000 57.190 653.145 58.235 ;
		LAYER M4 ;
		RECT 0.000 69.305 653.145 70.300 ;
		LAYER M4 ;
		RECT 0.000 71.110 653.145 72.155 ;
		LAYER M4 ;
		RECT 0.000 72.485 653.145 73.565 ;
		LAYER M4 ;
		RECT 0.000 73.945 653.145 74.940 ;
		LAYER M4 ;
		RECT 0.000 66.470 653.145 67.515 ;
		LAYER M4 ;
		RECT 0.000 83.225 653.535 84.220 ;
		LAYER M4 ;
		RECT 0.000 77.125 653.535 78.205 ;
		LAYER M4 ;
		RECT 0.000 80.390 653.535 81.435 ;
		LAYER M4 ;
		RECT 0.000 81.765 653.535 82.845 ;
		LAYER M4 ;
		RECT 0.000 75.750 653.535 76.795 ;
		LAYER M4 ;
		RECT 0.000 15.430 653.145 16.475 ;
		LAYER M4 ;
		RECT 0.000 13.625 653.145 14.620 ;
		LAYER M4 ;
		RECT 0.000 8.985 653.145 9.980 ;
		LAYER M4 ;
		RECT 0.000 7.525 653.145 8.605 ;
		LAYER M4 ;
		RECT 0.000 10.790 653.145 11.835 ;
		LAYER M4 ;
		RECT 0.000 12.165 653.145 13.245 ;
		LAYER M4 ;
		RECT 0.000 29.350 653.145 30.395 ;
		LAYER M4 ;
		RECT 0.000 24.710 653.145 25.755 ;
		LAYER M4 ;
		RECT 0.000 22.905 653.145 23.900 ;
		LAYER M4 ;
		RECT 0.000 26.085 653.145 27.165 ;
		LAYER M4 ;
		RECT 0.000 27.545 653.145 28.540 ;
		LAYER M4 ;
		RECT 0.000 30.725 653.145 31.805 ;
		LAYER M4 ;
		RECT 0.000 32.185 653.145 33.180 ;
		LAYER M4 ;
		RECT 0.000 33.990 653.145 35.035 ;
		LAYER M4 ;
		RECT 0.000 35.365 653.145 36.445 ;
		LAYER M4 ;
		RECT 0.000 36.825 653.145 37.820 ;
		LAYER M4 ;
		RECT 0.000 49.285 653.145 50.365 ;
		LAYER M4 ;
		RECT 0.000 46.105 653.145 47.100 ;
		LAYER M4 ;
		RECT 0.000 47.910 653.145 48.955 ;
		LAYER M4 ;
		RECT 0.000 50.745 653.145 51.740 ;
		LAYER M4 ;
		RECT 0.000 16.805 653.145 17.885 ;
		LAYER M4 ;
		RECT 0.000 18.265 653.145 19.260 ;
		LAYER M4 ;
		RECT 0.000 20.070 653.145 21.115 ;
		LAYER M4 ;
		RECT 0.000 21.445 653.145 22.525 ;
		LAYER M4 ;
		RECT 0.000 38.630 653.145 39.675 ;
		LAYER M4 ;
		RECT 0.000 41.465 653.145 42.460 ;
		LAYER M4 ;
		RECT 0.000 43.270 653.145 44.315 ;
		LAYER M4 ;
		RECT 0.000 44.645 653.145 45.725 ;
		LAYER M4 ;
		RECT 0.000 40.005 653.145 41.085 ;
	END
	# End of OBS

END TS1N28HPCPHVTB16384X36M8SSO

END LIBRARY
