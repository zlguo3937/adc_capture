# Created by MC2 : Version 2012.02.00.d on 2024/05/13, 17:41:26

#*********************************************************************************************************************/
# Software       : TSMC MEMORY COMPILER tsn28hpcpd127spsram_2012.02.00.d.180a						*/
# Technology     : TSMC 28nm CMOS LOGIC High Performance Compact Mobile Computing Plus 1P10M HKMG CU_ELK 0.9V				*/
#  Memory Type    : TSMC 28nm High Performance Compact Mobile Computing Plus Single Port SRAM with d127 bit cell SVT periphery */
# Library Name   : ts1n28hpcpsvtb32768x36m16swso (user specify : TS1N28HPCPSVTB32768X36M16SWSO)				*/
# Library Version: 180a												*/
# Generated Time : 2024/05/13, 17:41:17										*/
#*********************************************************************************************************************/
#															*/
# STATEMENT OF USE													*/
#															*/
# This information contains confidential and proprietary information of TSMC.					*/
# No part of this information may be reproduced, transmitted, transcribed,						*/
# stored in a retrieval system, or translated into any human or computer						*/
# language, in any form or by any means, electronic, mechanical, magnetic,						*/
# optical, chemical, manual, or otherwise, without the prior written permission					*/
# of TSMC. This information was prepared for informational purpose and is for					*/
# use by TSMC's customers only. TSMC reserves the right to make changes in the					*/
# information at any time and without notice.									*/
#															*/
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS1N28HPCPSVTB32768X36M16SWSO
	CLASS BLOCK ;
	FOREIGN TS1N28HPCPSVTB32768X36M16SWSO 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 654.735 BY 353.410 ;
	SYMMETRY X Y ;
	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 179.190 654.735 179.340 ;
			LAYER M1 ;
			RECT 654.555 179.190 654.735 179.340 ;
			LAYER M3 ;
			RECT 654.555 179.190 654.735 179.340 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[0]

	PIN A[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 169.330 654.735 169.480 ;
			LAYER M3 ;
			RECT 654.555 169.330 654.735 169.480 ;
			LAYER M2 ;
			RECT 654.555 169.330 654.735 169.480 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[10]

	PIN A[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 168.940 654.735 169.090 ;
			LAYER M2 ;
			RECT 654.555 168.940 654.735 169.090 ;
			LAYER M1 ;
			RECT 654.555 168.940 654.735 169.090 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[11]

	PIN A[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 181.630 654.735 181.780 ;
			LAYER M1 ;
			RECT 654.555 181.630 654.735 181.780 ;
			LAYER M2 ;
			RECT 654.555 181.630 654.735 181.780 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[12]

	PIN A[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 181.240 654.735 181.390 ;
			LAYER M2 ;
			RECT 654.555 181.240 654.735 181.390 ;
			LAYER M3 ;
			RECT 654.555 181.240 654.735 181.390 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[13]

	PIN A[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 179.580 654.735 179.730 ;
			LAYER M2 ;
			RECT 654.555 179.580 654.735 179.730 ;
			LAYER M1 ;
			RECT 654.555 179.580 654.735 179.730 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[14]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 177.530 654.735 177.680 ;
			LAYER M3 ;
			RECT 654.555 177.530 654.735 177.680 ;
			LAYER M2 ;
			RECT 654.555 177.530 654.735 177.680 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 177.140 654.735 177.290 ;
			LAYER M1 ;
			RECT 654.555 177.140 654.735 177.290 ;
			LAYER M3 ;
			RECT 654.555 177.140 654.735 177.290 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 167.280 654.735 167.430 ;
			LAYER M3 ;
			RECT 654.555 167.280 654.735 167.430 ;
			LAYER M2 ;
			RECT 654.555 167.280 654.735 167.430 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 173.040 654.735 173.190 ;
			LAYER M3 ;
			RECT 654.555 173.040 654.735 173.190 ;
			LAYER M1 ;
			RECT 654.555 173.040 654.735 173.190 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 171.380 654.735 171.530 ;
			LAYER M1 ;
			RECT 654.555 171.380 654.735 171.530 ;
			LAYER M2 ;
			RECT 654.555 171.380 654.735 171.530 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 170.990 654.735 171.140 ;
			LAYER M1 ;
			RECT 654.555 170.990 654.735 171.140 ;
			LAYER M2 ;
			RECT 654.555 170.990 654.735 171.140 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 175.480 654.735 175.630 ;
			LAYER M2 ;
			RECT 654.555 175.480 654.735 175.630 ;
			LAYER M3 ;
			RECT 654.555 175.480 654.735 175.630 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 175.090 654.735 175.240 ;
			LAYER M1 ;
			RECT 654.555 175.090 654.735 175.240 ;
			LAYER M2 ;
			RECT 654.555 175.090 654.735 175.240 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 173.430 654.735 173.580 ;
			LAYER M3 ;
			RECT 654.555 173.430 654.735 173.580 ;
			LAYER M1 ;
			RECT 654.555 173.430 654.735 173.580 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483700 LAYER M2 ;
		ANTENNAMAXAREACAR 18.165000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.065000 LAYER M3 ;
	END A[9]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 7.025 654.735 7.175 ;
			LAYER M2 ;
			RECT 654.555 7.025 654.735 7.175 ;
			LAYER M3 ;
			RECT 654.555 7.025 654.735 7.175 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 99.825 654.735 99.975 ;
			LAYER M1 ;
			RECT 654.555 99.825 654.735 99.975 ;
			LAYER M3 ;
			RECT 654.555 99.825 654.735 99.975 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 109.105 654.735 109.255 ;
			LAYER M1 ;
			RECT 654.555 109.105 654.735 109.255 ;
			LAYER M3 ;
			RECT 654.555 109.105 654.735 109.255 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 118.385 654.735 118.535 ;
			LAYER M1 ;
			RECT 654.555 118.385 654.735 118.535 ;
			LAYER M3 ;
			RECT 654.555 118.385 654.735 118.535 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 127.665 654.735 127.815 ;
			LAYER M3 ;
			RECT 654.555 127.665 654.735 127.815 ;
			LAYER M1 ;
			RECT 654.555 127.665 654.735 127.815 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 136.945 654.735 137.095 ;
			LAYER M3 ;
			RECT 654.555 136.945 654.735 137.095 ;
			LAYER M2 ;
			RECT 654.555 136.945 654.735 137.095 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 146.225 654.735 146.375 ;
			LAYER M3 ;
			RECT 654.555 146.225 654.735 146.375 ;
			LAYER M2 ;
			RECT 654.555 146.225 654.735 146.375 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 155.505 654.735 155.655 ;
			LAYER M3 ;
			RECT 654.555 155.505 654.735 155.655 ;
			LAYER M1 ;
			RECT 654.555 155.505 654.735 155.655 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 160.145 654.735 160.295 ;
			LAYER M1 ;
			RECT 654.555 160.145 654.735 160.295 ;
			LAYER M3 ;
			RECT 654.555 160.145 654.735 160.295 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 193.505 654.735 193.655 ;
			LAYER M3 ;
			RECT 654.555 193.505 654.735 193.655 ;
			LAYER M2 ;
			RECT 654.555 193.505 654.735 193.655 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 200.465 654.735 200.615 ;
			LAYER M1 ;
			RECT 654.555 200.465 654.735 200.615 ;
			LAYER M2 ;
			RECT 654.555 200.465 654.735 200.615 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 16.305 654.735 16.455 ;
			LAYER M2 ;
			RECT 654.555 16.305 654.735 16.455 ;
			LAYER M1 ;
			RECT 654.555 16.305 654.735 16.455 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 209.745 654.735 209.895 ;
			LAYER M2 ;
			RECT 654.555 209.745 654.735 209.895 ;
			LAYER M1 ;
			RECT 654.555 209.745 654.735 209.895 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 219.025 654.735 219.175 ;
			LAYER M1 ;
			RECT 654.555 219.025 654.735 219.175 ;
			LAYER M3 ;
			RECT 654.555 219.025 654.735 219.175 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 228.305 654.735 228.455 ;
			LAYER M3 ;
			RECT 654.555 228.305 654.735 228.455 ;
			LAYER M2 ;
			RECT 654.555 228.305 654.735 228.455 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 237.585 654.735 237.735 ;
			LAYER M3 ;
			RECT 654.555 237.585 654.735 237.735 ;
			LAYER M2 ;
			RECT 654.555 237.585 654.735 237.735 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 246.865 654.735 247.015 ;
			LAYER M3 ;
			RECT 654.555 246.865 654.735 247.015 ;
			LAYER M2 ;
			RECT 654.555 246.865 654.735 247.015 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 256.145 654.735 256.295 ;
			LAYER M3 ;
			RECT 654.555 256.145 654.735 256.295 ;
			LAYER M2 ;
			RECT 654.555 256.145 654.735 256.295 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 265.425 654.735 265.575 ;
			LAYER M1 ;
			RECT 654.555 265.425 654.735 265.575 ;
			LAYER M3 ;
			RECT 654.555 265.425 654.735 265.575 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 274.705 654.735 274.855 ;
			LAYER M1 ;
			RECT 654.555 274.705 654.735 274.855 ;
			LAYER M2 ;
			RECT 654.555 274.705 654.735 274.855 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 283.985 654.735 284.135 ;
			LAYER M3 ;
			RECT 654.555 283.985 654.735 284.135 ;
			LAYER M1 ;
			RECT 654.555 283.985 654.735 284.135 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 293.265 654.735 293.415 ;
			LAYER M3 ;
			RECT 654.555 293.265 654.735 293.415 ;
			LAYER M1 ;
			RECT 654.555 293.265 654.735 293.415 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 25.585 654.735 25.735 ;
			LAYER M2 ;
			RECT 654.555 25.585 654.735 25.735 ;
			LAYER M3 ;
			RECT 654.555 25.585 654.735 25.735 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 302.545 654.735 302.695 ;
			LAYER M3 ;
			RECT 654.555 302.545 654.735 302.695 ;
			LAYER M1 ;
			RECT 654.555 302.545 654.735 302.695 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 311.825 654.735 311.975 ;
			LAYER M2 ;
			RECT 654.555 311.825 654.735 311.975 ;
			LAYER M3 ;
			RECT 654.555 311.825 654.735 311.975 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[31]

	PIN BWEB[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 321.105 654.735 321.255 ;
			LAYER M1 ;
			RECT 654.555 321.105 654.735 321.255 ;
			LAYER M2 ;
			RECT 654.555 321.105 654.735 321.255 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[32]

	PIN BWEB[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 330.385 654.735 330.535 ;
			LAYER M2 ;
			RECT 654.555 330.385 654.735 330.535 ;
			LAYER M3 ;
			RECT 654.555 330.385 654.735 330.535 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[33]

	PIN BWEB[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 339.665 654.735 339.815 ;
			LAYER M1 ;
			RECT 654.555 339.665 654.735 339.815 ;
			LAYER M3 ;
			RECT 654.555 339.665 654.735 339.815 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[34]

	PIN BWEB[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 348.945 654.735 349.095 ;
			LAYER M2 ;
			RECT 654.555 348.945 654.735 349.095 ;
			LAYER M1 ;
			RECT 654.555 348.945 654.735 349.095 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[35]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 34.865 654.735 35.015 ;
			LAYER M3 ;
			RECT 654.555 34.865 654.735 35.015 ;
			LAYER M2 ;
			RECT 654.555 34.865 654.735 35.015 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 44.145 654.735 44.295 ;
			LAYER M2 ;
			RECT 654.555 44.145 654.735 44.295 ;
			LAYER M3 ;
			RECT 654.555 44.145 654.735 44.295 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 53.425 654.735 53.575 ;
			LAYER M2 ;
			RECT 654.555 53.425 654.735 53.575 ;
			LAYER M3 ;
			RECT 654.555 53.425 654.735 53.575 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 62.705 654.735 62.855 ;
			LAYER M2 ;
			RECT 654.555 62.705 654.735 62.855 ;
			LAYER M3 ;
			RECT 654.555 62.705 654.735 62.855 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 71.985 654.735 72.135 ;
			LAYER M2 ;
			RECT 654.555 71.985 654.735 72.135 ;
			LAYER M3 ;
			RECT 654.555 71.985 654.735 72.135 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 81.265 654.735 81.415 ;
			LAYER M1 ;
			RECT 654.555 81.265 654.735 81.415 ;
			LAYER M3 ;
			RECT 654.555 81.265 654.735 81.415 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 90.545 654.735 90.695 ;
			LAYER M1 ;
			RECT 654.555 90.545 654.735 90.695 ;
			LAYER M2 ;
			RECT 654.555 90.545 654.735 90.695 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.484400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.705000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.605000 LAYER M3 ;
	END BWEB[9]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 183.290 654.735 183.440 ;
			LAYER M2 ;
			RECT 654.555 183.290 654.735 183.440 ;
			LAYER M1 ;
			RECT 654.555 183.290 654.735 183.440 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.115300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.228300 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.515900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.249900 LAYER M2 ;
		ANTENNAMAXAREACAR 10.191100 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.732500 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 11.091100 LAYER M3 ;
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 183.920 654.735 184.070 ;
			LAYER M1 ;
			RECT 654.555 183.920 654.735 184.070 ;
			LAYER M2 ;
			RECT 654.555 183.920 654.735 184.070 ;
		END
		ANTENNAGATEAREA 2.013900 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 3.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 5.372500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.331500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA1 ;
		ANTENNAGATEAREA 2.013900 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 2.694600 LAYER M2 ;
		ANTENNAMAXAREACAR 33.912400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.292500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.097200 LAYER VIA2 ;
		ANTENNAGATEAREA 2.013900 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 2.754400 LAYER M3 ;
		ANTENNAMAXAREACAR 35.107800 LAYER M3 ;
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 6.635 654.735 6.785 ;
			LAYER M3 ;
			RECT 654.555 6.635 654.735 6.785 ;
			LAYER M2 ;
			RECT 654.555 6.635 654.735 6.785 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[0]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 99.435 654.735 99.585 ;
			LAYER M2 ;
			RECT 654.555 99.435 654.735 99.585 ;
			LAYER M1 ;
			RECT 654.555 99.435 654.735 99.585 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 108.715 654.735 108.865 ;
			LAYER M3 ;
			RECT 654.555 108.715 654.735 108.865 ;
			LAYER M1 ;
			RECT 654.555 108.715 654.735 108.865 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 117.995 654.735 118.145 ;
			LAYER M3 ;
			RECT 654.555 117.995 654.735 118.145 ;
			LAYER M1 ;
			RECT 654.555 117.995 654.735 118.145 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 127.275 654.735 127.425 ;
			LAYER M1 ;
			RECT 654.555 127.275 654.735 127.425 ;
			LAYER M3 ;
			RECT 654.555 127.275 654.735 127.425 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 136.555 654.735 136.705 ;
			LAYER M1 ;
			RECT 654.555 136.555 654.735 136.705 ;
			LAYER M3 ;
			RECT 654.555 136.555 654.735 136.705 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 145.835 654.735 145.985 ;
			LAYER M2 ;
			RECT 654.555 145.835 654.735 145.985 ;
			LAYER M1 ;
			RECT 654.555 145.835 654.735 145.985 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 155.115 654.735 155.265 ;
			LAYER M1 ;
			RECT 654.555 155.115 654.735 155.265 ;
			LAYER M3 ;
			RECT 654.555 155.115 654.735 155.265 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 159.755 654.735 159.905 ;
			LAYER M2 ;
			RECT 654.555 159.755 654.735 159.905 ;
			LAYER M3 ;
			RECT 654.555 159.755 654.735 159.905 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 193.115 654.735 193.265 ;
			LAYER M1 ;
			RECT 654.555 193.115 654.735 193.265 ;
			LAYER M2 ;
			RECT 654.555 193.115 654.735 193.265 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 200.075 654.735 200.225 ;
			LAYER M1 ;
			RECT 654.555 200.075 654.735 200.225 ;
			LAYER M3 ;
			RECT 654.555 200.075 654.735 200.225 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[19]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 15.915 654.735 16.065 ;
			LAYER M2 ;
			RECT 654.555 15.915 654.735 16.065 ;
			LAYER M1 ;
			RECT 654.555 15.915 654.735 16.065 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[1]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 209.355 654.735 209.505 ;
			LAYER M3 ;
			RECT 654.555 209.355 654.735 209.505 ;
			LAYER M2 ;
			RECT 654.555 209.355 654.735 209.505 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 218.635 654.735 218.785 ;
			LAYER M3 ;
			RECT 654.555 218.635 654.735 218.785 ;
			LAYER M1 ;
			RECT 654.555 218.635 654.735 218.785 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 227.915 654.735 228.065 ;
			LAYER M2 ;
			RECT 654.555 227.915 654.735 228.065 ;
			LAYER M3 ;
			RECT 654.555 227.915 654.735 228.065 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 237.195 654.735 237.345 ;
			LAYER M2 ;
			RECT 654.555 237.195 654.735 237.345 ;
			LAYER M3 ;
			RECT 654.555 237.195 654.735 237.345 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 246.475 654.735 246.625 ;
			LAYER M1 ;
			RECT 654.555 246.475 654.735 246.625 ;
			LAYER M2 ;
			RECT 654.555 246.475 654.735 246.625 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 255.755 654.735 255.905 ;
			LAYER M3 ;
			RECT 654.555 255.755 654.735 255.905 ;
			LAYER M1 ;
			RECT 654.555 255.755 654.735 255.905 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 265.035 654.735 265.185 ;
			LAYER M1 ;
			RECT 654.555 265.035 654.735 265.185 ;
			LAYER M2 ;
			RECT 654.555 265.035 654.735 265.185 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 274.315 654.735 274.465 ;
			LAYER M1 ;
			RECT 654.555 274.315 654.735 274.465 ;
			LAYER M2 ;
			RECT 654.555 274.315 654.735 274.465 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 283.595 654.735 283.745 ;
			LAYER M1 ;
			RECT 654.555 283.595 654.735 283.745 ;
			LAYER M2 ;
			RECT 654.555 283.595 654.735 283.745 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 292.875 654.735 293.025 ;
			LAYER M2 ;
			RECT 654.555 292.875 654.735 293.025 ;
			LAYER M1 ;
			RECT 654.555 292.875 654.735 293.025 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[29]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 25.195 654.735 25.345 ;
			LAYER M1 ;
			RECT 654.555 25.195 654.735 25.345 ;
			LAYER M2 ;
			RECT 654.555 25.195 654.735 25.345 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[2]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 302.155 654.735 302.305 ;
			LAYER M1 ;
			RECT 654.555 302.155 654.735 302.305 ;
			LAYER M3 ;
			RECT 654.555 302.155 654.735 302.305 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 311.435 654.735 311.585 ;
			LAYER M1 ;
			RECT 654.555 311.435 654.735 311.585 ;
			LAYER M3 ;
			RECT 654.555 311.435 654.735 311.585 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[31]

	PIN D[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 320.715 654.735 320.865 ;
			LAYER M2 ;
			RECT 654.555 320.715 654.735 320.865 ;
			LAYER M3 ;
			RECT 654.555 320.715 654.735 320.865 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[32]

	PIN D[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 329.995 654.735 330.145 ;
			LAYER M1 ;
			RECT 654.555 329.995 654.735 330.145 ;
			LAYER M2 ;
			RECT 654.555 329.995 654.735 330.145 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[33]

	PIN D[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 339.275 654.735 339.425 ;
			LAYER M3 ;
			RECT 654.555 339.275 654.735 339.425 ;
			LAYER M1 ;
			RECT 654.555 339.275 654.735 339.425 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[34]

	PIN D[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 348.555 654.735 348.705 ;
			LAYER M3 ;
			RECT 654.555 348.555 654.735 348.705 ;
			LAYER M2 ;
			RECT 654.555 348.555 654.735 348.705 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[35]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 34.475 654.735 34.625 ;
			LAYER M3 ;
			RECT 654.555 34.475 654.735 34.625 ;
			LAYER M2 ;
			RECT 654.555 34.475 654.735 34.625 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 43.755 654.735 43.905 ;
			LAYER M2 ;
			RECT 654.555 43.755 654.735 43.905 ;
			LAYER M1 ;
			RECT 654.555 43.755 654.735 43.905 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 53.035 654.735 53.185 ;
			LAYER M3 ;
			RECT 654.555 53.035 654.735 53.185 ;
			LAYER M1 ;
			RECT 654.555 53.035 654.735 53.185 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 62.315 654.735 62.465 ;
			LAYER M3 ;
			RECT 654.555 62.315 654.735 62.465 ;
			LAYER M1 ;
			RECT 654.555 62.315 654.735 62.465 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 71.595 654.735 71.745 ;
			LAYER M2 ;
			RECT 654.555 71.595 654.735 71.745 ;
			LAYER M3 ;
			RECT 654.555 71.595 654.735 71.745 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 80.875 654.735 81.025 ;
			LAYER M1 ;
			RECT 654.555 80.875 654.735 81.025 ;
			LAYER M2 ;
			RECT 654.555 80.875 654.735 81.025 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 90.155 654.735 90.305 ;
			LAYER M1 ;
			RECT 654.555 90.155 654.735 90.305 ;
			LAYER M2 ;
			RECT 654.555 90.155 654.735 90.305 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.125300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.560000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.481400 LAYER M2 ;
		ANTENNAMAXAREACAR 18.608300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 19.508300 LAYER M3 ;
	END D[9]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 7.645 654.735 7.795 ;
			LAYER M3 ;
			RECT 654.555 7.645 654.735 7.795 ;
			LAYER M1 ;
			RECT 654.555 7.645 654.735 7.795 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[0]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 100.445 654.735 100.595 ;
			LAYER M2 ;
			RECT 654.555 100.445 654.735 100.595 ;
			LAYER M3 ;
			RECT 654.555 100.445 654.735 100.595 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 109.725 654.735 109.875 ;
			LAYER M2 ;
			RECT 654.555 109.725 654.735 109.875 ;
			LAYER M3 ;
			RECT 654.555 109.725 654.735 109.875 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 119.005 654.735 119.155 ;
			LAYER M2 ;
			RECT 654.555 119.005 654.735 119.155 ;
			LAYER M1 ;
			RECT 654.555 119.005 654.735 119.155 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 128.285 654.735 128.435 ;
			LAYER M3 ;
			RECT 654.555 128.285 654.735 128.435 ;
			LAYER M2 ;
			RECT 654.555 128.285 654.735 128.435 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 137.565 654.735 137.715 ;
			LAYER M2 ;
			RECT 654.555 137.565 654.735 137.715 ;
			LAYER M3 ;
			RECT 654.555 137.565 654.735 137.715 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 146.845 654.735 146.995 ;
			LAYER M3 ;
			RECT 654.555 146.845 654.735 146.995 ;
			LAYER M1 ;
			RECT 654.555 146.845 654.735 146.995 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 156.125 654.735 156.275 ;
			LAYER M2 ;
			RECT 654.555 156.125 654.735 156.275 ;
			LAYER M1 ;
			RECT 654.555 156.125 654.735 156.275 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 160.765 654.735 160.915 ;
			LAYER M3 ;
			RECT 654.555 160.765 654.735 160.915 ;
			LAYER M1 ;
			RECT 654.555 160.765 654.735 160.915 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 194.125 654.735 194.275 ;
			LAYER M1 ;
			RECT 654.555 194.125 654.735 194.275 ;
			LAYER M3 ;
			RECT 654.555 194.125 654.735 194.275 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 201.085 654.735 201.235 ;
			LAYER M3 ;
			RECT 654.555 201.085 654.735 201.235 ;
			LAYER M2 ;
			RECT 654.555 201.085 654.735 201.235 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[19]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 16.925 654.735 17.075 ;
			LAYER M1 ;
			RECT 654.555 16.925 654.735 17.075 ;
			LAYER M2 ;
			RECT 654.555 16.925 654.735 17.075 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[1]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 210.365 654.735 210.515 ;
			LAYER M1 ;
			RECT 654.555 210.365 654.735 210.515 ;
			LAYER M3 ;
			RECT 654.555 210.365 654.735 210.515 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 219.645 654.735 219.795 ;
			LAYER M2 ;
			RECT 654.555 219.645 654.735 219.795 ;
			LAYER M1 ;
			RECT 654.555 219.645 654.735 219.795 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 228.925 654.735 229.075 ;
			LAYER M2 ;
			RECT 654.555 228.925 654.735 229.075 ;
			LAYER M3 ;
			RECT 654.555 228.925 654.735 229.075 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 238.205 654.735 238.355 ;
			LAYER M3 ;
			RECT 654.555 238.205 654.735 238.355 ;
			LAYER M2 ;
			RECT 654.555 238.205 654.735 238.355 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 247.485 654.735 247.635 ;
			LAYER M1 ;
			RECT 654.555 247.485 654.735 247.635 ;
			LAYER M3 ;
			RECT 654.555 247.485 654.735 247.635 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 256.765 654.735 256.915 ;
			LAYER M2 ;
			RECT 654.555 256.765 654.735 256.915 ;
			LAYER M3 ;
			RECT 654.555 256.765 654.735 256.915 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 266.045 654.735 266.195 ;
			LAYER M1 ;
			RECT 654.555 266.045 654.735 266.195 ;
			LAYER M2 ;
			RECT 654.555 266.045 654.735 266.195 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 275.325 654.735 275.475 ;
			LAYER M2 ;
			RECT 654.555 275.325 654.735 275.475 ;
			LAYER M3 ;
			RECT 654.555 275.325 654.735 275.475 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 284.605 654.735 284.755 ;
			LAYER M1 ;
			RECT 654.555 284.605 654.735 284.755 ;
			LAYER M2 ;
			RECT 654.555 284.605 654.735 284.755 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 293.885 654.735 294.035 ;
			LAYER M2 ;
			RECT 654.555 293.885 654.735 294.035 ;
			LAYER M1 ;
			RECT 654.555 293.885 654.735 294.035 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[29]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 26.205 654.735 26.355 ;
			LAYER M1 ;
			RECT 654.555 26.205 654.735 26.355 ;
			LAYER M3 ;
			RECT 654.555 26.205 654.735 26.355 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[2]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 303.165 654.735 303.315 ;
			LAYER M3 ;
			RECT 654.555 303.165 654.735 303.315 ;
			LAYER M1 ;
			RECT 654.555 303.165 654.735 303.315 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 312.445 654.735 312.595 ;
			LAYER M1 ;
			RECT 654.555 312.445 654.735 312.595 ;
			LAYER M3 ;
			RECT 654.555 312.445 654.735 312.595 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[31]

	PIN Q[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 321.725 654.735 321.875 ;
			LAYER M1 ;
			RECT 654.555 321.725 654.735 321.875 ;
			LAYER M3 ;
			RECT 654.555 321.725 654.735 321.875 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[32]

	PIN Q[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 331.005 654.735 331.155 ;
			LAYER M2 ;
			RECT 654.555 331.005 654.735 331.155 ;
			LAYER M3 ;
			RECT 654.555 331.005 654.735 331.155 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[33]

	PIN Q[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 340.285 654.735 340.435 ;
			LAYER M2 ;
			RECT 654.555 340.285 654.735 340.435 ;
			LAYER M3 ;
			RECT 654.555 340.285 654.735 340.435 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[34]

	PIN Q[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 349.565 654.735 349.715 ;
			LAYER M1 ;
			RECT 654.555 349.565 654.735 349.715 ;
			LAYER M2 ;
			RECT 654.555 349.565 654.735 349.715 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[35]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 35.485 654.735 35.635 ;
			LAYER M2 ;
			RECT 654.555 35.485 654.735 35.635 ;
			LAYER M3 ;
			RECT 654.555 35.485 654.735 35.635 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 44.765 654.735 44.915 ;
			LAYER M1 ;
			RECT 654.555 44.765 654.735 44.915 ;
			LAYER M2 ;
			RECT 654.555 44.765 654.735 44.915 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 54.045 654.735 54.195 ;
			LAYER M3 ;
			RECT 654.555 54.045 654.735 54.195 ;
			LAYER M1 ;
			RECT 654.555 54.045 654.735 54.195 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 63.325 654.735 63.475 ;
			LAYER M2 ;
			RECT 654.555 63.325 654.735 63.475 ;
			LAYER M3 ;
			RECT 654.555 63.325 654.735 63.475 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 72.605 654.735 72.755 ;
			LAYER M3 ;
			RECT 654.555 72.605 654.735 72.755 ;
			LAYER M2 ;
			RECT 654.555 72.605 654.735 72.755 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 81.885 654.735 82.035 ;
			LAYER M2 ;
			RECT 654.555 81.885 654.735 82.035 ;
			LAYER M3 ;
			RECT 654.555 81.885 654.735 82.035 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 654.555 91.165 654.735 91.315 ;
			LAYER M3 ;
			RECT 654.555 91.165 654.735 91.315 ;
			LAYER M2 ;
			RECT 654.555 91.165 654.735 91.315 ;
		END
		ANTENNADIFFAREA 0.163000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.265500 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.163000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.154000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.163000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.176700 LAYER M3 ;
	END Q[9]

	PIN SD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 654.555 164.665 654.735 164.815 ;
			LAYER M2 ;
			RECT 654.555 164.665 654.735 164.815 ;
			LAYER M1 ;
			RECT 654.555 164.665 654.735 164.815 ;
		END
		ANTENNAGATEAREA 0.051000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.839700 LAYER M1 ;
		ANTENNAMAXAREACAR 9.087800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.585600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.051000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.499900 LAYER M2 ;
		ANTENNAMAXAREACAR 48.990700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.878400 LAYER VIA2 ;
		ANTENNAGATEAREA 0.051000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.590600 LAYER M3 ;
		ANTENNAMAXAREACAR 48.990700 LAYER M3 ;
	END SD

	PIN SLP
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 165.380 654.735 165.530 ;
			LAYER M1 ;
			RECT 654.555 165.380 654.735 165.530 ;
			LAYER M3 ;
			RECT 654.555 165.380 654.735 165.530 ;
		END
		ANTENNAGATEAREA 0.027000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.172400 LAYER M1 ;
		ANTENNAMAXAREACAR 8.260000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.433300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.027000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.269000 LAYER M2 ;
		ANTENNAMAXAREACAR 48.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.027000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.564300 LAYER M3 ;
		ANTENNAMAXAREACAR 48.814800 LAYER M3 ;
	END SLP

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.000 4.875 654.345 5.205 ;
			LAYER M4 ;
			RECT 0.000 14.155 654.345 14.485 ;
			LAYER M4 ;
			RECT 0.000 23.435 654.345 23.765 ;
			LAYER M4 ;
			RECT 0.000 32.715 654.345 33.045 ;
			LAYER M4 ;
			RECT 0.000 41.995 654.345 42.325 ;
			LAYER M4 ;
			RECT 0.000 51.275 654.345 51.605 ;
			LAYER M4 ;
			RECT 0.000 60.555 654.345 60.885 ;
			LAYER M4 ;
			RECT 0.000 69.835 654.345 70.165 ;
			LAYER M4 ;
			RECT 0.000 79.115 654.345 79.445 ;
			LAYER M4 ;
			RECT 0.000 88.395 654.345 88.725 ;
			LAYER M4 ;
			RECT 0.000 97.675 654.345 98.005 ;
			LAYER M4 ;
			RECT 0.000 106.955 654.345 107.285 ;
			LAYER M4 ;
			RECT 0.000 116.235 654.345 116.565 ;
			LAYER M4 ;
			RECT 0.000 125.515 654.345 125.845 ;
			LAYER M4 ;
			RECT 0.000 134.795 654.345 135.125 ;
			LAYER M4 ;
			RECT 0.000 144.075 654.345 144.405 ;
			LAYER M4 ;
			RECT 0.000 153.355 654.345 153.685 ;
			LAYER M4 ;
			RECT 0.000 162.635 654.735 162.965 ;
			LAYER M4 ;
			RECT 0.000 175.275 654.735 175.845 ;
			LAYER M4 ;
			RECT 0.000 175.975 654.735 176.545 ;
			LAYER M4 ;
			RECT 0.000 182.955 654.735 183.525 ;
			LAYER M4 ;
			RECT 0.000 189.035 654.735 189.365 ;
			LAYER M4 ;
			RECT 0.000 198.315 654.345 198.645 ;
			LAYER M4 ;
			RECT 0.000 207.595 654.345 207.925 ;
			LAYER M4 ;
			RECT 0.000 216.875 654.345 217.205 ;
			LAYER M4 ;
			RECT 0.000 226.155 654.345 226.485 ;
			LAYER M4 ;
			RECT 0.000 235.435 654.345 235.765 ;
			LAYER M4 ;
			RECT 0.000 244.715 654.345 245.045 ;
			LAYER M4 ;
			RECT 0.000 253.995 654.345 254.325 ;
			LAYER M4 ;
			RECT 0.000 263.275 654.345 263.605 ;
			LAYER M4 ;
			RECT 0.000 272.555 654.345 272.885 ;
			LAYER M4 ;
			RECT 0.000 281.835 654.345 282.165 ;
			LAYER M4 ;
			RECT 0.000 291.115 654.345 291.445 ;
			LAYER M4 ;
			RECT 0.000 300.395 654.345 300.725 ;
			LAYER M4 ;
			RECT 0.000 309.675 654.345 310.005 ;
			LAYER M4 ;
			RECT 0.000 318.955 654.345 319.285 ;
			LAYER M4 ;
			RECT 0.000 328.235 654.345 328.565 ;
			LAYER M4 ;
			RECT 0.000 337.515 654.345 337.845 ;
			LAYER M4 ;
			RECT 0.000 346.795 654.345 347.125 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.000 6.285 654.345 6.665 ;
			LAYER M4 ;
			RECT 0.000 15.565 654.345 15.945 ;
			LAYER M4 ;
			RECT 0.000 24.845 654.345 25.225 ;
			LAYER M4 ;
			RECT 0.000 34.125 654.345 34.505 ;
			LAYER M4 ;
			RECT 0.000 43.405 654.345 43.785 ;
			LAYER M4 ;
			RECT 0.000 52.685 654.345 53.065 ;
			LAYER M4 ;
			RECT 0.000 61.965 654.345 62.345 ;
			LAYER M4 ;
			RECT 0.000 71.245 654.345 71.625 ;
			LAYER M4 ;
			RECT 0.000 80.525 654.345 80.905 ;
			LAYER M4 ;
			RECT 0.000 89.805 654.345 90.185 ;
			LAYER M4 ;
			RECT 0.000 99.085 654.345 99.465 ;
			LAYER M4 ;
			RECT 0.000 108.365 654.345 108.745 ;
			LAYER M4 ;
			RECT 0.000 117.645 654.345 118.025 ;
			LAYER M4 ;
			RECT 0.000 126.925 654.345 127.305 ;
			LAYER M4 ;
			RECT 0.000 136.205 654.345 136.585 ;
			LAYER M4 ;
			RECT 0.000 145.485 654.345 145.865 ;
			LAYER M4 ;
			RECT 0.000 154.765 654.345 155.145 ;
			LAYER M4 ;
			RECT 0.000 164.045 654.735 164.425 ;
			LAYER M4 ;
			RECT 0.000 173.875 654.735 174.445 ;
			LAYER M4 ;
			RECT 0.000 174.575 654.735 175.145 ;
			LAYER M4 ;
			RECT 0.000 176.905 654.735 177.475 ;
			LAYER M4 ;
			RECT 0.000 190.445 654.735 190.825 ;
			LAYER M4 ;
			RECT 0.000 199.725 654.345 200.105 ;
			LAYER M4 ;
			RECT 0.000 209.005 654.345 209.385 ;
			LAYER M4 ;
			RECT 0.000 218.285 654.345 218.665 ;
			LAYER M4 ;
			RECT 0.000 227.565 654.345 227.945 ;
			LAYER M4 ;
			RECT 0.000 236.845 654.345 237.225 ;
			LAYER M4 ;
			RECT 0.000 246.125 654.345 246.505 ;
			LAYER M4 ;
			RECT 0.000 255.405 654.345 255.785 ;
			LAYER M4 ;
			RECT 0.000 264.685 654.345 265.065 ;
			LAYER M4 ;
			RECT 0.000 273.965 654.345 274.345 ;
			LAYER M4 ;
			RECT 0.000 283.245 654.345 283.625 ;
			LAYER M4 ;
			RECT 0.000 292.525 654.345 292.905 ;
			LAYER M4 ;
			RECT 0.000 301.805 654.345 302.185 ;
			LAYER M4 ;
			RECT 0.000 311.085 654.345 311.465 ;
			LAYER M4 ;
			RECT 0.000 320.365 654.345 320.745 ;
			LAYER M4 ;
			RECT 0.000 329.645 654.345 330.025 ;
			LAYER M4 ;
			RECT 0.000 338.925 654.345 339.305 ;
			LAYER M4 ;
			RECT 0.000 348.205 654.345 348.585 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 654.555 166.890 654.735 167.040 ;
			LAYER M3 ;
			RECT 654.555 166.890 654.735 167.040 ;
			LAYER M1 ;
			RECT 654.555 166.890 654.735 167.040 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.109700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.041700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.445400 LAYER M2 ;
		ANTENNAMAXAREACAR 16.888300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.500000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 17.788300 LAYER M3 ;
	END WEB

	OBS
		# Promoted blockages
		LAYER M1 ;
		RECT 654.555 303.375 654.735 311.375 ;
		LAYER M1 ;
		RECT 654.555 312.655 654.735 320.655 ;
		LAYER M3 ;
		RECT 654.555 312.675 654.735 320.635 ;
		LAYER M2 ;
		RECT 654.555 303.395 654.735 311.355 ;
		LAYER M3 ;
		RECT 654.555 303.395 654.735 311.355 ;
		LAYER VIA3 ;
		RECT 654.555 303.395 654.735 311.355 ;
		LAYER M3 ;
		RECT 654.555 321.335 654.735 321.645 ;
		LAYER VIA3 ;
		RECT 654.555 321.335 654.735 321.645 ;
		LAYER VIA3 ;
		RECT 654.555 312.675 654.735 320.635 ;
		LAYER M3 ;
		RECT 654.555 320.945 654.735 321.025 ;
		LAYER M1 ;
		RECT 654.555 320.925 654.735 321.045 ;
		LAYER VIA3 ;
		RECT 654.555 320.945 654.735 321.025 ;
		LAYER M2 ;
		RECT 654.555 321.335 654.735 321.645 ;
		LAYER M1 ;
		RECT 654.555 321.315 654.735 321.665 ;
		LAYER M2 ;
		RECT 654.555 320.945 654.735 321.025 ;
		LAYER M2 ;
		RECT 654.555 312.675 654.735 320.635 ;
		LAYER M2 ;
		RECT 654.555 302.775 654.735 303.085 ;
		LAYER M1 ;
		RECT 654.555 302.365 654.735 302.485 ;
		LAYER M2 ;
		RECT 654.555 294.115 654.735 302.075 ;
		LAYER VIA3 ;
		RECT 654.555 294.115 654.735 302.075 ;
		LAYER M3 ;
		RECT 654.555 294.115 654.735 302.075 ;
		LAYER M1 ;
		RECT 654.555 294.095 654.735 302.095 ;
		LAYER VIA3 ;
		RECT 654.555 284.835 654.735 292.795 ;
		LAYER M1 ;
		RECT 654.555 284.815 654.735 292.815 ;
		LAYER M2 ;
		RECT 654.555 293.105 654.735 293.185 ;
		LAYER M3 ;
		RECT 654.555 293.105 654.735 293.185 ;
		LAYER M3 ;
		RECT 654.555 284.835 654.735 292.795 ;
		LAYER VIA3 ;
		RECT 654.555 283.825 654.735 283.905 ;
		LAYER M2 ;
		RECT 654.555 284.215 654.735 284.525 ;
		LAYER M3 ;
		RECT 654.555 284.215 654.735 284.525 ;
		LAYER M1 ;
		RECT 654.555 275.535 654.735 283.535 ;
		LAYER M1 ;
		RECT 654.555 293.085 654.735 293.205 ;
		LAYER M2 ;
		RECT 654.555 293.495 654.735 293.805 ;
		LAYER M3 ;
		RECT 654.555 275.555 654.735 283.515 ;
		LAYER VIA3 ;
		RECT 654.555 275.555 654.735 283.515 ;
		LAYER M1 ;
		RECT 654.555 302.755 654.735 303.105 ;
		LAYER VIA3 ;
		RECT 654.555 302.385 654.735 302.465 ;
		LAYER M2 ;
		RECT 654.555 302.385 654.735 302.465 ;
		LAYER M3 ;
		RECT 654.555 302.385 654.735 302.465 ;
		LAYER VIA3 ;
		RECT 654.555 302.775 654.735 303.085 ;
		LAYER M1 ;
		RECT 654.555 274.915 654.735 275.265 ;
		LAYER M2 ;
		RECT 654.555 274.935 654.735 275.245 ;
		LAYER M3 ;
		RECT 654.555 274.935 654.735 275.245 ;
		LAYER M2 ;
		RECT 654.555 274.545 654.735 274.625 ;
		LAYER M3 ;
		RECT 654.555 274.545 654.735 274.625 ;
		LAYER M3 ;
		RECT 654.555 293.495 654.735 293.805 ;
		LAYER M1 ;
		RECT 654.555 293.475 654.735 293.825 ;
		LAYER M1 ;
		RECT 654.555 274.525 654.735 274.645 ;
		LAYER M2 ;
		RECT 654.555 330.225 654.735 330.305 ;
		LAYER M2 ;
		RECT 654.555 331.235 654.735 339.195 ;
		LAYER M3 ;
		RECT 654.555 331.235 654.735 339.195 ;
		LAYER M3 ;
		RECT 654.555 330.615 654.735 330.925 ;
		LAYER M1 ;
		RECT 654.555 330.595 654.735 330.945 ;
		LAYER VIA3 ;
		RECT 654.555 330.225 654.735 330.305 ;
		LAYER M2 ;
		RECT 654.555 339.895 654.735 340.205 ;
		LAYER VIA3 ;
		RECT 654.555 339.895 654.735 340.205 ;
		LAYER M3 ;
		RECT 654.555 339.895 654.735 340.205 ;
		LAYER M2 ;
		RECT 654.555 339.505 654.735 339.585 ;
		LAYER VIA3 ;
		RECT 654.555 339.505 654.735 339.585 ;
		LAYER M3 ;
		RECT 654.555 339.505 654.735 339.585 ;
		LAYER M3 ;
		RECT 654.555 330.225 654.735 330.305 ;
		LAYER M1 ;
		RECT 654.555 339.875 654.735 340.225 ;
		LAYER M1 ;
		RECT 654.555 339.485 654.735 339.605 ;
		LAYER M1 ;
		RECT 654.555 331.215 654.735 339.215 ;
		LAYER M2 ;
		RECT 654.555 340.515 654.735 348.475 ;
		LAYER M1 ;
		RECT 654.555 340.495 654.735 348.495 ;
		LAYER M2 ;
		RECT 654.555 348.785 654.735 348.865 ;
		LAYER M3 ;
		RECT 654.555 348.785 654.735 348.865 ;
		LAYER VIA3 ;
		RECT 654.555 348.785 654.735 348.865 ;
		LAYER M3 ;
		RECT 654.555 340.515 654.735 348.475 ;
		LAYER VIA3 ;
		RECT 654.555 340.515 654.735 348.475 ;
		LAYER M1 ;
		RECT 654.555 348.765 654.735 348.885 ;
		LAYER M1 ;
		RECT 654.555 330.205 654.735 330.325 ;
		LAYER VIA3 ;
		RECT 654.555 330.615 654.735 330.925 ;
		LAYER M2 ;
		RECT 654.555 330.615 654.735 330.925 ;
		LAYER VIA3 ;
		RECT 654.555 331.235 654.735 339.195 ;
		LAYER M1 ;
		RECT 654.555 349.155 654.735 349.505 ;
		LAYER M2 ;
		RECT 654.555 349.175 654.735 349.485 ;
		LAYER M3 ;
		RECT 654.555 349.175 654.735 349.485 ;
		LAYER VIA3 ;
		RECT 654.555 349.175 654.735 349.485 ;
		LAYER M1 ;
		RECT 654.555 349.775 654.735 353.410 ;
		LAYER M2 ;
		RECT 654.555 349.795 654.735 353.410 ;
		LAYER M3 ;
		RECT 654.555 349.795 654.735 353.410 ;
		LAYER VIA3 ;
		RECT 654.555 349.795 654.735 353.410 ;
		LAYER M2 ;
		RECT 654.555 321.955 654.735 329.915 ;
		LAYER M3 ;
		RECT 654.555 321.955 654.735 329.915 ;
		LAYER VIA3 ;
		RECT 654.555 321.955 654.735 329.915 ;
		LAYER M1 ;
		RECT 654.555 321.935 654.735 329.935 ;
		LAYER M2 ;
		RECT 654.555 53.265 654.735 53.345 ;
		LAYER M2 ;
		RECT 654.555 53.655 654.735 53.965 ;
		LAYER M3 ;
		RECT 654.555 53.655 654.735 53.965 ;
		LAYER M2 ;
		RECT 654.555 63.555 654.735 71.515 ;
		LAYER M3 ;
		RECT 654.555 53.265 654.735 53.345 ;
		LAYER VIA3 ;
		RECT 654.555 53.265 654.735 53.345 ;
		LAYER M3 ;
		RECT 654.555 63.555 654.735 71.515 ;
		LAYER M2 ;
		RECT 654.555 7.875 654.735 15.835 ;
		LAYER M2 ;
		RECT 654.555 7.255 654.735 7.565 ;
		LAYER M1 ;
		RECT 654.555 7.235 654.735 7.585 ;
		LAYER M1 ;
		RECT 654.555 6.845 654.735 6.965 ;
		LAYER M3 ;
		RECT 654.555 7.255 654.735 7.565 ;
		LAYER M3 ;
		RECT 654.555 7.875 654.735 15.835 ;
		LAYER M2 ;
		RECT 654.555 16.535 654.735 16.845 ;
		LAYER M1 ;
		RECT 654.555 16.515 654.735 16.865 ;
		LAYER M3 ;
		RECT 654.555 16.535 654.735 16.845 ;
		LAYER VIA3 ;
		RECT 654.555 16.145 654.735 16.225 ;
		LAYER M3 ;
		RECT 654.555 82.115 654.735 90.075 ;
		LAYER M2 ;
		RECT 654.555 90.775 654.735 91.085 ;
		LAYER M3 ;
		RECT 654.555 90.775 654.735 91.085 ;
		LAYER VIA3 ;
		RECT 654.555 90.775 654.735 91.085 ;
		LAYER M1 ;
		RECT 654.555 100.655 654.735 108.655 ;
		LAYER M2 ;
		RECT 654.555 100.675 654.735 108.635 ;
		LAYER M2 ;
		RECT 654.555 100.055 654.735 100.365 ;
		LAYER M1 ;
		RECT 654.555 100.035 654.735 100.385 ;
		LAYER M2 ;
		RECT 654.555 91.395 654.735 99.355 ;
		LAYER M2 ;
		RECT 654.555 108.945 654.735 109.025 ;
		LAYER M1 ;
		RECT 654.555 108.925 654.735 109.045 ;
		LAYER M1 ;
		RECT 654.555 109.935 654.735 117.935 ;
		LAYER VIA3 ;
		RECT 654.555 118.225 654.735 118.305 ;
		LAYER M2 ;
		RECT 654.555 118.225 654.735 118.305 ;
		LAYER M3 ;
		RECT 654.555 118.225 654.735 118.305 ;
		LAYER M2 ;
		RECT 654.555 109.955 654.735 117.915 ;
		LAYER VIA3 ;
		RECT 654.555 109.955 654.735 117.915 ;
		LAYER M3 ;
		RECT 654.555 109.955 654.735 117.915 ;
		LAYER M2 ;
		RECT 654.555 109.335 654.735 109.645 ;
		LAYER VIA3 ;
		RECT 654.555 109.335 654.735 109.645 ;
		LAYER M3 ;
		RECT 654.555 109.335 654.735 109.645 ;
		LAYER M1 ;
		RECT 654.555 109.315 654.735 109.665 ;
		LAYER M3 ;
		RECT 654.555 81.495 654.735 81.805 ;
		LAYER M2 ;
		RECT 654.555 128.515 654.735 136.475 ;
		LAYER M3 ;
		RECT 654.555 128.515 654.735 136.475 ;
		LAYER M1 ;
		RECT 654.555 118.205 654.735 118.325 ;
		LAYER M2 ;
		RECT 654.555 137.795 654.735 145.755 ;
		LAYER M2 ;
		RECT 654.555 146.455 654.735 146.765 ;
		LAYER M3 ;
		RECT 654.555 146.455 654.735 146.765 ;
		LAYER VIA3 ;
		RECT 654.555 159.985 654.735 160.065 ;
		LAYER M3 ;
		RECT 654.555 156.355 654.735 159.675 ;
		LAYER M3 ;
		RECT 654.555 155.735 654.735 156.045 ;
		LAYER M1 ;
		RECT 654.555 155.715 654.735 156.065 ;
		LAYER VIA3 ;
		RECT 654.555 160.375 654.735 160.685 ;
		LAYER M3 ;
		RECT 654.555 160.375 654.735 160.685 ;
		LAYER M2 ;
		RECT 654.555 159.985 654.735 160.065 ;
		LAYER M3 ;
		RECT 654.555 159.985 654.735 160.065 ;
		LAYER M2 ;
		RECT 654.555 90.385 654.735 90.465 ;
		LAYER M3 ;
		RECT 654.555 90.385 654.735 90.465 ;
		LAYER M2 ;
		RECT 654.555 72.215 654.735 72.525 ;
		LAYER M3 ;
		RECT 654.555 72.215 654.735 72.525 ;
		LAYER M1 ;
		RECT 654.555 82.095 654.735 90.095 ;
		LAYER VIA3 ;
		RECT 654.555 160.995 654.735 164.585 ;
		LAYER M1 ;
		RECT 654.555 147.055 654.735 155.055 ;
		LAYER M2 ;
		RECT 654.555 147.075 654.735 155.035 ;
		LAYER M1 ;
		RECT 654.555 160.355 654.735 160.705 ;
		LAYER M2 ;
		RECT 654.555 155.345 654.735 155.425 ;
		LAYER M1 ;
		RECT 654.555 155.325 654.735 155.445 ;
		LAYER M4 ;
		RECT 389.275 6.665 406.505 7.195 ;
		LAYER M4 ;
		RECT 389.275 29.110 406.505 30.990 ;
		LAYER M4 ;
		RECT 389.275 26.900 406.505 28.945 ;
		LAYER M4 ;
		RECT 389.275 25.225 406.505 25.755 ;
		LAYER M4 ;
		RECT 389.275 4.735 406.505 4.875 ;
		LAYER M4 ;
		RECT 389.275 32.575 406.505 32.715 ;
		LAYER M4 ;
		RECT 389.275 34.505 406.505 35.035 ;
		LAYER M4 ;
		RECT 389.275 36.180 406.505 38.225 ;
		LAYER M4 ;
		RECT 389.275 38.390 406.505 40.270 ;
		LAYER M4 ;
		RECT 71.735 6.665 88.965 7.195 ;
		LAYER M4 ;
		RECT 247.735 6.665 389.275 7.160 ;
		LAYER M4 ;
		RECT 389.275 15.945 406.505 16.475 ;
		LAYER M4 ;
		RECT 71.735 8.340 88.965 10.385 ;
		LAYER M4 ;
		RECT 88.965 6.665 230.505 7.160 ;
		LAYER M4 ;
		RECT 389.275 8.340 406.505 10.385 ;
		LAYER M4 ;
		RECT 389.275 14.015 406.505 14.155 ;
		LAYER M4 ;
		RECT 389.275 17.620 406.505 19.665 ;
		LAYER M4 ;
		RECT 389.275 19.830 406.505 21.710 ;
		LAYER M4 ;
		RECT 389.275 10.550 406.505 12.430 ;
		LAYER M4 ;
		RECT 389.275 88.255 406.505 88.395 ;
		LAYER M4 ;
		RECT 389.275 56.950 406.505 58.830 ;
		LAYER M4 ;
		RECT 389.275 53.065 406.505 53.595 ;
		LAYER M4 ;
		RECT 389.275 84.790 406.505 86.670 ;
		LAYER M4 ;
		RECT 389.275 82.580 406.505 84.625 ;
		LAYER M4 ;
		RECT 389.275 80.905 406.505 81.435 ;
		LAYER M4 ;
		RECT 389.275 73.300 406.505 75.345 ;
		LAYER M4 ;
		RECT 0.000 32.575 1.365 32.715 ;
		LAYER M4 ;
		RECT 0.000 33.045 654.345 34.125 ;
		LAYER M4 ;
		RECT 0.000 23.765 654.345 24.845 ;
		LAYER M4 ;
		RECT 0.000 51.605 654.345 52.685 ;
		LAYER M4 ;
		RECT 0.000 23.295 1.365 23.435 ;
		LAYER M4 ;
		RECT 0.000 4.735 1.365 4.875 ;
		LAYER M4 ;
		RECT 0.000 5.205 654.345 6.285 ;
		LAYER M4 ;
		RECT 0.000 41.855 1.365 41.995 ;
		LAYER M4 ;
		RECT 0.000 34.505 71.735 35.000 ;
		LAYER M4 ;
		RECT 71.735 51.135 88.965 51.275 ;
		LAYER M4 ;
		RECT 71.735 1.270 88.965 3.150 ;
		LAYER M4 ;
		RECT 71.735 330.025 88.965 330.555 ;
		LAYER M4 ;
		RECT 71.735 333.910 88.965 335.790 ;
		LAYER M4 ;
		RECT 71.735 337.375 88.965 337.515 ;
		LAYER M1 ;
		RECT 654.555 0.000 654.735 6.575 ;
		LAYER M2 ;
		RECT 654.555 0.000 654.735 6.555 ;
		LAYER M3 ;
		RECT 654.555 0.000 654.735 6.555 ;
		LAYER M4 ;
		RECT 0.000 162.965 654.735 164.045 ;
		LAYER VIA3 ;
		RECT 654.555 0.000 654.735 6.555 ;
		LAYER M4 ;
		RECT 388.675 183.525 654.735 185.060 ;
		LAYER M4 ;
		RECT 0.000 189.365 654.735 190.445 ;
		LAYER M4 ;
		RECT 0.000 177.475 654.735 182.955 ;
		LAYER M4 ;
		RECT 0.000 168.055 654.735 173.875 ;
		LAYER M4 ;
		RECT 230.505 331.700 247.735 333.745 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 654.735 353.410 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 654.735 353.410 ;
		LAYER M2 ;
		RECT 654.555 82.115 654.735 90.075 ;
		LAYER VIA3 ;
		RECT 654.555 82.115 654.735 90.075 ;
		LAYER M1 ;
		RECT 654.555 91.375 654.735 99.375 ;
		LAYER M3 ;
		RECT 654.555 72.835 654.735 80.795 ;
		LAYER M3 ;
		RECT 654.555 100.675 654.735 108.635 ;
		LAYER M3 ;
		RECT 654.555 108.945 654.735 109.025 ;
		LAYER VIA3 ;
		RECT 654.555 100.675 654.735 108.635 ;
		LAYER VIA3 ;
		RECT 654.555 108.945 654.735 109.025 ;
		LAYER M2 ;
		RECT 654.555 99.665 654.735 99.745 ;
		LAYER M1 ;
		RECT 654.555 99.645 654.735 99.765 ;
		LAYER M3 ;
		RECT 654.555 100.055 654.735 100.365 ;
		LAYER M3 ;
		RECT 654.555 99.665 654.735 99.745 ;
		LAYER VIA3 ;
		RECT 654.555 99.665 654.735 99.745 ;
		LAYER VIA3 ;
		RECT 654.555 100.055 654.735 100.365 ;
		LAYER M1 ;
		RECT 654.555 90.755 654.735 91.105 ;
		LAYER VIA3 ;
		RECT 654.555 90.385 654.735 90.465 ;
		LAYER M1 ;
		RECT 654.555 90.365 654.735 90.485 ;
		LAYER VIA3 ;
		RECT 654.555 91.395 654.735 99.355 ;
		LAYER M3 ;
		RECT 654.555 91.395 654.735 99.355 ;
		LAYER M2 ;
		RECT 654.555 81.495 654.735 81.805 ;
		LAYER M2 ;
		RECT 654.555 62.545 654.735 62.625 ;
		LAYER M3 ;
		RECT 654.555 62.545 654.735 62.625 ;
		LAYER VIA3 ;
		RECT 654.555 62.545 654.735 62.625 ;
		LAYER M1 ;
		RECT 654.555 81.085 654.735 81.205 ;
		LAYER M3 ;
		RECT 654.555 71.825 654.735 71.905 ;
		LAYER VIA3 ;
		RECT 654.555 71.825 654.735 71.905 ;
		LAYER VIA3 ;
		RECT 654.555 81.105 654.735 81.185 ;
		LAYER M1 ;
		RECT 654.555 72.195 654.735 72.545 ;
		LAYER M2 ;
		RECT 654.555 71.825 654.735 71.905 ;
		LAYER M2 ;
		RECT 654.555 81.105 654.735 81.185 ;
		LAYER M3 ;
		RECT 654.555 81.105 654.735 81.185 ;
		LAYER VIA3 ;
		RECT 654.555 63.555 654.735 71.515 ;
		LAYER M1 ;
		RECT 654.555 71.805 654.735 71.925 ;
		LAYER M1 ;
		RECT 654.555 81.475 654.735 81.825 ;
		LAYER M2 ;
		RECT 654.555 62.935 654.735 63.245 ;
		LAYER M3 ;
		RECT 654.555 62.935 654.735 63.245 ;
		LAYER VIA3 ;
		RECT 654.555 62.935 654.735 63.245 ;
		LAYER VIA3 ;
		RECT 654.555 81.495 654.735 81.805 ;
		LAYER M1 ;
		RECT 654.555 63.535 654.735 71.535 ;
		LAYER M2 ;
		RECT 654.555 72.835 654.735 80.795 ;
		LAYER VIA3 ;
		RECT 654.555 72.835 654.735 80.795 ;
		LAYER M1 ;
		RECT 654.555 72.815 654.735 80.815 ;
		LAYER VIA3 ;
		RECT 654.555 72.215 654.735 72.525 ;
		LAYER M1 ;
		RECT 654.555 137.155 654.735 137.505 ;
		LAYER M2 ;
		RECT 654.555 136.785 654.735 136.865 ;
		LAYER M3 ;
		RECT 654.555 136.785 654.735 136.865 ;
		LAYER VIA3 ;
		RECT 654.555 136.785 654.735 136.865 ;
		LAYER M2 ;
		RECT 654.555 137.175 654.735 137.485 ;
		LAYER M3 ;
		RECT 654.555 137.175 654.735 137.485 ;
		LAYER VIA3 ;
		RECT 654.555 137.175 654.735 137.485 ;
		LAYER VIA3 ;
		RECT 654.555 146.455 654.735 146.765 ;
		LAYER M1 ;
		RECT 654.555 136.765 654.735 136.885 ;
		LAYER VIA3 ;
		RECT 654.555 128.515 654.735 136.475 ;
		LAYER M1 ;
		RECT 654.555 128.495 654.735 136.495 ;
		LAYER M1 ;
		RECT 654.555 146.435 654.735 146.785 ;
		LAYER M2 ;
		RECT 654.555 119.235 654.735 127.195 ;
		LAYER M3 ;
		RECT 654.555 119.235 654.735 127.195 ;
		LAYER M2 ;
		RECT 654.555 118.615 654.735 118.925 ;
		LAYER VIA3 ;
		RECT 654.555 147.075 654.735 155.035 ;
		LAYER M1 ;
		RECT 654.555 137.775 654.735 145.775 ;
		LAYER M3 ;
		RECT 654.555 137.795 654.735 145.755 ;
		LAYER VIA3 ;
		RECT 654.555 137.795 654.735 145.755 ;
		LAYER M2 ;
		RECT 654.555 146.065 654.735 146.145 ;
		LAYER M3 ;
		RECT 654.555 146.065 654.735 146.145 ;
		LAYER VIA3 ;
		RECT 654.555 146.065 654.735 146.145 ;
		LAYER M1 ;
		RECT 654.555 146.045 654.735 146.165 ;
		LAYER M3 ;
		RECT 654.555 147.075 654.735 155.035 ;
		LAYER M1 ;
		RECT 654.555 164.875 654.735 165.320 ;
		LAYER M3 ;
		RECT 654.555 160.995 654.735 164.585 ;
		LAYER M2 ;
		RECT 654.555 160.995 654.735 164.585 ;
		LAYER M1 ;
		RECT 654.555 160.975 654.735 164.605 ;
		LAYER M2 ;
		RECT 654.555 127.895 654.735 128.205 ;
		LAYER M3 ;
		RECT 654.555 127.895 654.735 128.205 ;
		LAYER M1 ;
		RECT 654.555 127.485 654.735 127.605 ;
		LAYER M1 ;
		RECT 654.555 127.875 654.735 128.225 ;
		LAYER M2 ;
		RECT 654.555 127.505 654.735 127.585 ;
		LAYER M3 ;
		RECT 654.555 127.505 654.735 127.585 ;
		LAYER VIA3 ;
		RECT 654.555 127.505 654.735 127.585 ;
		LAYER VIA3 ;
		RECT 654.555 127.895 654.735 128.205 ;
		LAYER M3 ;
		RECT 654.555 118.615 654.735 118.925 ;
		LAYER VIA3 ;
		RECT 654.555 118.615 654.735 118.925 ;
		LAYER M1 ;
		RECT 654.555 118.595 654.735 118.945 ;
		LAYER VIA3 ;
		RECT 654.555 119.235 654.735 127.195 ;
		LAYER M1 ;
		RECT 654.555 119.215 654.735 127.215 ;
		LAYER M3 ;
		RECT 654.555 44.995 654.735 52.955 ;
		LAYER M2 ;
		RECT 654.555 35.715 654.735 43.675 ;
		LAYER VIA3 ;
		RECT 654.555 35.715 654.735 43.675 ;
		LAYER M2 ;
		RECT 654.555 54.275 654.735 62.235 ;
		LAYER VIA3 ;
		RECT 654.555 53.655 654.735 53.965 ;
		LAYER M1 ;
		RECT 654.555 53.245 654.735 53.365 ;
		LAYER M1 ;
		RECT 654.555 43.965 654.735 44.085 ;
		LAYER M2 ;
		RECT 654.555 44.375 654.735 44.685 ;
		LAYER M3 ;
		RECT 654.555 44.375 654.735 44.685 ;
		LAYER M1 ;
		RECT 654.555 44.355 654.735 44.705 ;
		LAYER VIA3 ;
		RECT 654.555 44.375 654.735 44.685 ;
		LAYER VIA3 ;
		RECT 654.555 44.995 654.735 52.955 ;
		LAYER M1 ;
		RECT 654.555 25.795 654.735 26.145 ;
		LAYER VIA3 ;
		RECT 654.555 25.425 654.735 25.505 ;
		LAYER M2 ;
		RECT 654.555 43.985 654.735 44.065 ;
		LAYER M3 ;
		RECT 654.555 43.985 654.735 44.065 ;
		LAYER VIA3 ;
		RECT 654.555 43.985 654.735 44.065 ;
		LAYER M1 ;
		RECT 654.555 26.415 654.735 34.415 ;
		LAYER M2 ;
		RECT 654.555 26.435 654.735 34.395 ;
		LAYER VIA3 ;
		RECT 654.555 26.435 654.735 34.395 ;
		LAYER M2 ;
		RECT 654.555 25.815 654.735 26.125 ;
		LAYER M3 ;
		RECT 654.555 25.815 654.735 26.125 ;
		LAYER M2 ;
		RECT 654.555 35.095 654.735 35.405 ;
		LAYER M3 ;
		RECT 654.555 35.095 654.735 35.405 ;
		LAYER VIA3 ;
		RECT 654.555 25.815 654.735 26.125 ;
		LAYER M1 ;
		RECT 654.555 35.695 654.735 43.695 ;
		LAYER VIA3 ;
		RECT 654.555 35.095 654.735 35.405 ;
		LAYER M1 ;
		RECT 654.555 35.075 654.735 35.425 ;
		LAYER M3 ;
		RECT 654.555 35.715 654.735 43.675 ;
		LAYER M1 ;
		RECT 654.555 17.135 654.735 25.135 ;
		LAYER M2 ;
		RECT 654.555 17.155 654.735 25.115 ;
		LAYER M2 ;
		RECT 654.555 25.425 654.735 25.505 ;
		LAYER M3 ;
		RECT 654.555 25.425 654.735 25.505 ;
		LAYER M3 ;
		RECT 654.555 17.155 654.735 25.115 ;
		LAYER VIA3 ;
		RECT 654.555 17.155 654.735 25.115 ;
		LAYER M3 ;
		RECT 654.555 34.705 654.735 34.785 ;
		LAYER M2 ;
		RECT 654.555 34.705 654.735 34.785 ;
		LAYER VIA3 ;
		RECT 654.555 34.705 654.735 34.785 ;
		LAYER M1 ;
		RECT 654.555 34.685 654.735 34.805 ;
		LAYER M1 ;
		RECT 654.555 169.540 654.735 170.930 ;
		LAYER M1 ;
		RECT 654.555 167.100 654.735 167.220 ;
		LAYER M1 ;
		RECT 654.555 165.590 654.735 166.830 ;
		LAYER VIA3 ;
		RECT 654.555 164.895 654.735 165.300 ;
		LAYER M1 ;
		RECT 654.555 167.490 654.735 168.880 ;
		LAYER M1 ;
		RECT 654.555 169.150 654.735 169.270 ;
		LAYER M3 ;
		RECT 654.555 169.170 654.735 169.250 ;
		LAYER M3 ;
		RECT 654.555 167.510 654.735 168.860 ;
		LAYER VIA3 ;
		RECT 654.555 167.510 654.735 168.860 ;
		LAYER VIA3 ;
		RECT 654.555 169.170 654.735 169.250 ;
		LAYER M2 ;
		RECT 654.555 167.120 654.735 167.200 ;
		LAYER M3 ;
		RECT 654.555 167.120 654.735 167.200 ;
		LAYER M2 ;
		RECT 654.555 165.610 654.735 166.810 ;
		LAYER VIA3 ;
		RECT 654.555 167.120 654.735 167.200 ;
		LAYER M3 ;
		RECT 654.555 165.610 654.735 166.810 ;
		LAYER VIA3 ;
		RECT 654.555 165.610 654.735 166.810 ;
		LAYER M2 ;
		RECT 654.555 155.735 654.735 156.045 ;
		LAYER VIA3 ;
		RECT 654.555 155.735 654.735 156.045 ;
		LAYER M3 ;
		RECT 654.555 155.345 654.735 155.425 ;
		LAYER VIA3 ;
		RECT 654.555 156.355 654.735 159.675 ;
		LAYER VIA3 ;
		RECT 654.555 155.345 654.735 155.425 ;
		LAYER M1 ;
		RECT 654.555 183.500 654.735 183.860 ;
		LAYER M2 ;
		RECT 654.555 194.355 654.735 199.995 ;
		LAYER M1 ;
		RECT 654.555 194.335 654.735 200.015 ;
		LAYER M2 ;
		RECT 654.555 201.315 654.735 209.275 ;
		LAYER M1 ;
		RECT 654.555 200.285 654.735 200.405 ;
		LAYER M3 ;
		RECT 654.555 229.155 654.735 237.115 ;
		LAYER M1 ;
		RECT 654.555 219.855 654.735 227.855 ;
		LAYER M1 ;
		RECT 654.555 219.235 654.735 219.585 ;
		LAYER M2 ;
		RECT 654.555 229.155 654.735 237.115 ;
		LAYER M1 ;
		RECT 654.555 229.135 654.735 237.135 ;
		LAYER M2 ;
		RECT 654.555 228.535 654.735 228.845 ;
		LAYER M3 ;
		RECT 654.555 228.535 654.735 228.845 ;
		LAYER VIA3 ;
		RECT 654.555 228.535 654.735 228.845 ;
		LAYER VIA3 ;
		RECT 654.555 229.155 654.735 237.115 ;
		LAYER M2 ;
		RECT 654.555 228.145 654.735 228.225 ;
		LAYER M3 ;
		RECT 654.555 228.145 654.735 228.225 ;
		LAYER VIA3 ;
		RECT 654.555 228.145 654.735 228.225 ;
		LAYER M1 ;
		RECT 654.555 228.125 654.735 228.245 ;
		LAYER M1 ;
		RECT 654.555 228.515 654.735 228.865 ;
		LAYER M2 ;
		RECT 654.555 219.875 654.735 227.835 ;
		LAYER M3 ;
		RECT 654.555 219.875 654.735 227.835 ;
		LAYER VIA3 ;
		RECT 654.555 219.875 654.735 227.835 ;
		LAYER M1 ;
		RECT 654.555 201.295 654.735 209.295 ;
		LAYER M2 ;
		RECT 654.555 209.585 654.735 209.665 ;
		LAYER M3 ;
		RECT 654.555 209.585 654.735 209.665 ;
		LAYER VIA3 ;
		RECT 654.555 209.585 654.735 209.665 ;
		LAYER M3 ;
		RECT 654.555 201.315 654.735 209.275 ;
		LAYER VIA3 ;
		RECT 654.555 201.315 654.735 209.275 ;
		LAYER M1 ;
		RECT 654.555 209.955 654.735 210.305 ;
		LAYER VIA3 ;
		RECT 654.555 209.975 654.735 210.285 ;
		LAYER M2 ;
		RECT 654.555 209.975 654.735 210.285 ;
		LAYER M3 ;
		RECT 654.555 209.975 654.735 210.285 ;
		LAYER M1 ;
		RECT 654.555 210.575 654.735 218.575 ;
		LAYER VIA3 ;
		RECT 654.555 210.595 654.735 218.555 ;
		LAYER M2 ;
		RECT 654.555 218.865 654.735 218.945 ;
		LAYER M3 ;
		RECT 654.555 218.865 654.735 218.945 ;
		LAYER VIA3 ;
		RECT 654.555 218.865 654.735 218.945 ;
		LAYER M1 ;
		RECT 654.555 218.845 654.735 218.965 ;
		LAYER M2 ;
		RECT 654.555 200.695 654.735 201.005 ;
		LAYER M3 ;
		RECT 654.555 200.695 654.735 201.005 ;
		LAYER M1 ;
		RECT 654.555 200.675 654.735 201.025 ;
		LAYER VIA3 ;
		RECT 654.555 200.695 654.735 201.005 ;
		LAYER M2 ;
		RECT 654.555 210.595 654.735 218.555 ;
		LAYER M3 ;
		RECT 654.555 210.595 654.735 218.555 ;
		LAYER M1 ;
		RECT 654.555 209.565 654.735 209.685 ;
		LAYER M2 ;
		RECT 654.555 219.255 654.735 219.565 ;
		LAYER M3 ;
		RECT 654.555 219.255 654.735 219.565 ;
		LAYER VIA3 ;
		RECT 654.555 219.255 654.735 219.565 ;
		LAYER M1 ;
		RECT 654.555 181.840 654.735 183.230 ;
		LAYER M3 ;
		RECT 654.555 183.520 654.735 183.840 ;
		LAYER VIA3 ;
		RECT 654.555 183.520 654.735 183.840 ;
		LAYER VIA3 ;
		RECT 654.555 184.150 654.735 193.035 ;
		LAYER VIA3 ;
		RECT 654.555 181.470 654.735 181.550 ;
		LAYER M2 ;
		RECT 654.555 181.860 654.735 183.210 ;
		LAYER M3 ;
		RECT 654.555 181.860 654.735 183.210 ;
		LAYER VIA3 ;
		RECT 654.555 181.860 654.735 183.210 ;
		LAYER M3 ;
		RECT 654.555 193.345 654.735 193.425 ;
		LAYER M2 ;
		RECT 654.555 200.305 654.735 200.385 ;
		LAYER M3 ;
		RECT 654.555 200.305 654.735 200.385 ;
		LAYER VIA3 ;
		RECT 654.555 193.345 654.735 193.425 ;
		LAYER VIA3 ;
		RECT 654.555 200.305 654.735 200.385 ;
		LAYER M3 ;
		RECT 654.555 193.735 654.735 194.045 ;
		LAYER VIA3 ;
		RECT 654.555 193.735 654.735 194.045 ;
		LAYER VIA3 ;
		RECT 654.555 194.355 654.735 199.995 ;
		LAYER M3 ;
		RECT 654.555 194.355 654.735 199.995 ;
		LAYER M1 ;
		RECT 654.555 173.640 654.735 175.030 ;
		LAYER M2 ;
		RECT 654.555 173.660 654.735 175.010 ;
		LAYER M3 ;
		RECT 654.555 173.660 654.735 175.010 ;
		LAYER VIA3 ;
		RECT 654.555 173.660 654.735 175.010 ;
		LAYER M1 ;
		RECT 654.555 175.300 654.735 175.420 ;
		LAYER M1 ;
		RECT 654.555 177.350 654.735 177.470 ;
		LAYER M2 ;
		RECT 654.555 177.370 654.735 177.450 ;
		LAYER VIA3 ;
		RECT 654.555 175.320 654.735 175.400 ;
		LAYER M3 ;
		RECT 654.555 177.370 654.735 177.450 ;
		LAYER VIA3 ;
		RECT 654.555 177.370 654.735 177.450 ;
		LAYER M2 ;
		RECT 654.555 175.320 654.735 175.400 ;
		LAYER M3 ;
		RECT 654.555 175.320 654.735 175.400 ;
		LAYER M2 ;
		RECT 654.555 177.760 654.735 179.110 ;
		LAYER M3 ;
		RECT 654.555 177.760 654.735 179.110 ;
		LAYER VIA3 ;
		RECT 654.555 177.760 654.735 179.110 ;
		LAYER M3 ;
		RECT 654.555 171.220 654.735 171.300 ;
		LAYER VIA3 ;
		RECT 654.555 171.220 654.735 171.300 ;
		LAYER M2 ;
		RECT 654.555 171.610 654.735 172.960 ;
		LAYER M3 ;
		RECT 654.555 171.610 654.735 172.960 ;
		LAYER M1 ;
		RECT 654.555 171.590 654.735 172.980 ;
		LAYER M1 ;
		RECT 654.555 177.740 654.735 179.130 ;
		LAYER M1 ;
		RECT 654.555 173.250 654.735 173.370 ;
		LAYER VIA3 ;
		RECT 654.555 171.610 654.735 172.960 ;
		LAYER M2 ;
		RECT 654.555 179.810 654.735 181.160 ;
		LAYER M3 ;
		RECT 654.555 179.810 654.735 181.160 ;
		LAYER VIA3 ;
		RECT 654.555 179.420 654.735 179.500 ;
		LAYER M2 ;
		RECT 654.555 175.710 654.735 177.060 ;
		LAYER M3 ;
		RECT 654.555 175.710 654.735 177.060 ;
		LAYER VIA3 ;
		RECT 654.555 175.710 654.735 177.060 ;
		LAYER M1 ;
		RECT 654.555 175.690 654.735 177.080 ;
		LAYER M2 ;
		RECT 654.555 183.520 654.735 183.840 ;
		LAYER M1 ;
		RECT 654.555 193.325 654.735 193.445 ;
		LAYER M1 ;
		RECT 654.555 193.715 654.735 194.065 ;
		LAYER M2 ;
		RECT 654.555 193.735 654.735 194.045 ;
		LAYER M2 ;
		RECT 654.555 256.375 654.735 256.685 ;
		LAYER M1 ;
		RECT 654.555 256.355 654.735 256.705 ;
		LAYER M2 ;
		RECT 654.555 256.995 654.735 264.955 ;
		LAYER M3 ;
		RECT 654.555 256.995 654.735 264.955 ;
		LAYER M3 ;
		RECT 654.555 256.375 654.735 256.685 ;
		LAYER VIA3 ;
		RECT 654.555 256.375 654.735 256.685 ;
		LAYER VIA3 ;
		RECT 654.555 256.995 654.735 264.955 ;
		LAYER M1 ;
		RECT 654.555 184.130 654.735 193.055 ;
		LAYER M2 ;
		RECT 654.555 184.150 654.735 193.035 ;
		LAYER M3 ;
		RECT 654.555 184.150 654.735 193.035 ;
		LAYER M2 ;
		RECT 654.555 193.345 654.735 193.425 ;
		LAYER M1 ;
		RECT 654.555 237.795 654.735 238.145 ;
		LAYER M2 ;
		RECT 654.555 265.265 654.735 265.345 ;
		LAYER M1 ;
		RECT 654.555 247.075 654.735 247.425 ;
		LAYER M3 ;
		RECT 654.555 265.265 654.735 265.345 ;
		LAYER VIA3 ;
		RECT 654.555 265.265 654.735 265.345 ;
		LAYER M1 ;
		RECT 654.555 256.975 654.735 264.975 ;
		LAYER M2 ;
		RECT 654.555 237.425 654.735 237.505 ;
		LAYER M3 ;
		RECT 654.555 265.655 654.735 265.965 ;
		LAYER VIA3 ;
		RECT 654.555 265.655 654.735 265.965 ;
		LAYER M1 ;
		RECT 654.555 265.245 654.735 265.365 ;
		LAYER M2 ;
		RECT 654.555 265.655 654.735 265.965 ;
		LAYER M2 ;
		RECT 654.555 171.220 654.735 171.300 ;
		LAYER M2 ;
		RECT 654.555 173.270 654.735 173.350 ;
		LAYER M3 ;
		RECT 654.555 173.270 654.735 173.350 ;
		LAYER VIA3 ;
		RECT 654.555 173.270 654.735 173.350 ;
		LAYER M2 ;
		RECT 654.555 169.560 654.735 170.910 ;
		LAYER M3 ;
		RECT 654.555 179.420 654.735 179.500 ;
		LAYER M1 ;
		RECT 654.555 179.400 654.735 179.520 ;
		LAYER M3 ;
		RECT 654.555 169.560 654.735 170.910 ;
		LAYER VIA3 ;
		RECT 654.555 169.560 654.735 170.910 ;
		LAYER M1 ;
		RECT 654.555 171.200 654.735 171.320 ;
		LAYER M1 ;
		RECT 654.555 179.790 654.735 181.180 ;
		LAYER M2 ;
		RECT 654.555 181.470 654.735 181.550 ;
		LAYER M1 ;
		RECT 654.555 181.450 654.735 181.570 ;
		LAYER M2 ;
		RECT 654.555 179.420 654.735 179.500 ;
		LAYER VIA3 ;
		RECT 654.555 179.810 654.735 181.160 ;
		LAYER M3 ;
		RECT 654.555 181.470 654.735 181.550 ;
		LAYER M2 ;
		RECT 654.555 238.435 654.735 246.395 ;
		LAYER M3 ;
		RECT 654.555 238.435 654.735 246.395 ;
		LAYER VIA3 ;
		RECT 654.555 238.435 654.735 246.395 ;
		LAYER M2 ;
		RECT 654.555 246.705 654.735 246.785 ;
		LAYER M3 ;
		RECT 654.555 237.425 654.735 237.505 ;
		LAYER M1 ;
		RECT 654.555 237.405 654.735 237.525 ;
		LAYER VIA3 ;
		RECT 654.555 246.705 654.735 246.785 ;
		LAYER M3 ;
		RECT 654.555 246.705 654.735 246.785 ;
		LAYER M1 ;
		RECT 654.555 246.685 654.735 246.805 ;
		LAYER M2 ;
		RECT 654.555 247.095 654.735 247.405 ;
		LAYER M3 ;
		RECT 654.555 247.095 654.735 247.405 ;
		LAYER VIA3 ;
		RECT 654.555 247.095 654.735 247.405 ;
		LAYER M2 ;
		RECT 654.555 255.985 654.735 256.065 ;
		LAYER M1 ;
		RECT 654.555 255.965 654.735 256.085 ;
		LAYER M2 ;
		RECT 654.555 247.715 654.735 255.675 ;
		LAYER VIA3 ;
		RECT 654.555 247.715 654.735 255.675 ;
		LAYER M3 ;
		RECT 654.555 237.815 654.735 238.125 ;
		LAYER M2 ;
		RECT 654.555 237.815 654.735 238.125 ;
		LAYER VIA3 ;
		RECT 654.555 237.815 654.735 238.125 ;
		LAYER VIA3 ;
		RECT 654.555 237.425 654.735 237.505 ;
		LAYER M3 ;
		RECT 654.555 255.985 654.735 256.065 ;
		LAYER VIA3 ;
		RECT 654.555 255.985 654.735 256.065 ;
		LAYER M3 ;
		RECT 654.555 247.715 654.735 255.675 ;
		LAYER M4 ;
		RECT 548.045 302.185 565.275 302.715 ;
		LAYER M4 ;
		RECT 548.045 300.255 565.275 300.395 ;
		LAYER M4 ;
		RECT 548.045 296.790 565.275 298.670 ;
		LAYER M4 ;
		RECT 548.045 294.580 565.275 296.625 ;
		LAYER M4 ;
		RECT 548.045 309.535 565.275 309.675 ;
		LAYER M4 ;
		RECT 548.045 313.140 565.275 315.185 ;
		LAYER M4 ;
		RECT 548.045 315.350 565.275 317.230 ;
		LAYER M4 ;
		RECT 548.045 318.815 565.275 318.955 ;
		LAYER M4 ;
		RECT 548.045 311.465 565.275 311.995 ;
		LAYER M4 ;
		RECT 548.045 226.015 565.275 226.155 ;
		LAYER M4 ;
		RECT 548.045 128.980 565.275 131.025 ;
		LAYER M4 ;
		RECT 548.045 127.305 565.275 127.835 ;
		LAYER M4 ;
		RECT 548.045 121.910 565.275 123.790 ;
		LAYER M4 ;
		RECT 548.045 125.375 565.275 125.515 ;
		LAYER M4 ;
		RECT 548.045 119.700 565.275 121.745 ;
		LAYER M4 ;
		RECT 548.045 118.025 565.275 118.555 ;
		LAYER M4 ;
		RECT 548.045 303.860 565.275 305.905 ;
		LAYER M4 ;
		RECT 548.045 292.905 565.275 293.435 ;
		LAYER M4 ;
		RECT 548.045 290.975 565.275 291.115 ;
		LAYER M4 ;
		RECT 548.045 287.510 565.275 289.390 ;
		LAYER M4 ;
		RECT 548.045 306.070 565.275 307.950 ;
		LAYER M4 ;
		RECT 548.045 285.300 565.275 287.345 ;
		LAYER M4 ;
		RECT 548.045 283.625 565.275 284.155 ;
		LAYER M4 ;
		RECT 548.045 227.945 565.275 228.475 ;
		LAYER M4 ;
		RECT 548.045 241.110 565.275 242.990 ;
		LAYER M4 ;
		RECT 548.045 218.665 565.275 219.195 ;
		LAYER M4 ;
		RECT 548.045 222.550 565.275 224.430 ;
		LAYER M4 ;
		RECT 548.045 231.830 565.275 233.710 ;
		LAYER M4 ;
		RECT 548.045 235.295 565.275 235.435 ;
		LAYER M4 ;
		RECT 548.045 229.620 565.275 231.665 ;
		LAYER M4 ;
		RECT 548.045 238.900 565.275 240.945 ;
		LAYER M4 ;
		RECT 548.045 237.225 565.275 237.755 ;
		LAYER M4 ;
		RECT 548.045 131.190 565.275 133.070 ;
		LAYER M4 ;
		RECT 548.045 201.780 565.275 203.825 ;
		LAYER M4 ;
		RECT 548.045 200.105 565.275 200.635 ;
		LAYER M4 ;
		RECT 548.045 10.550 565.275 12.430 ;
		LAYER M4 ;
		RECT 548.045 15.945 565.275 16.475 ;
		LAYER M4 ;
		RECT 548.045 17.620 565.275 19.665 ;
		LAYER M4 ;
		RECT 548.045 19.830 565.275 21.710 ;
		LAYER M4 ;
		RECT 548.045 14.015 565.275 14.155 ;
		LAYER M4 ;
		RECT 548.045 8.340 565.275 10.385 ;
		LAYER M4 ;
		RECT 548.045 101.140 565.275 103.185 ;
		LAYER M4 ;
		RECT 548.045 103.350 565.275 105.230 ;
		LAYER M4 ;
		RECT 548.045 106.815 565.275 106.955 ;
		LAYER M4 ;
		RECT 548.045 110.420 565.275 112.465 ;
		LAYER M4 ;
		RECT 548.045 112.630 565.275 114.510 ;
		LAYER M4 ;
		RECT 548.045 116.095 565.275 116.235 ;
		LAYER M4 ;
		RECT 548.045 99.465 565.275 99.995 ;
		LAYER M4 ;
		RECT 548.045 78.975 565.275 79.115 ;
		LAYER M4 ;
		RECT 548.045 71.625 565.275 72.155 ;
		LAYER M4 ;
		RECT 548.045 25.225 565.275 25.755 ;
		LAYER M4 ;
		RECT 548.045 23.295 565.275 23.435 ;
		LAYER M4 ;
		RECT 548.045 26.900 565.275 28.945 ;
		LAYER M4 ;
		RECT 548.045 29.110 565.275 30.990 ;
		LAYER M4 ;
		RECT 548.045 32.575 565.275 32.715 ;
		LAYER M4 ;
		RECT 548.045 36.180 565.275 38.225 ;
		LAYER M4 ;
		RECT 548.045 38.390 565.275 40.270 ;
		LAYER M4 ;
		RECT 548.045 41.855 565.275 41.995 ;
		LAYER M4 ;
		RECT 548.045 43.785 565.275 44.315 ;
		LAYER M4 ;
		RECT 548.045 34.505 565.275 35.035 ;
		LAYER M4 ;
		RECT 548.045 54.740 565.275 56.785 ;
		LAYER M4 ;
		RECT 548.045 56.950 565.275 58.830 ;
		LAYER M4 ;
		RECT 548.045 97.535 565.275 97.675 ;
		LAYER M4 ;
		RECT 548.045 66.230 565.275 68.110 ;
		LAYER M4 ;
		RECT 548.045 73.300 565.275 75.345 ;
		LAYER M4 ;
		RECT 548.045 94.070 565.275 95.950 ;
		LAYER M4 ;
		RECT 548.045 91.860 565.275 93.905 ;
		LAYER M4 ;
		RECT 548.045 60.415 565.275 60.555 ;
		LAYER M4 ;
		RECT 548.045 88.255 565.275 88.395 ;
		LAYER M4 ;
		RECT 548.045 82.580 565.275 84.625 ;
		LAYER M4 ;
		RECT 548.045 80.905 565.275 81.435 ;
		LAYER M4 ;
		RECT 548.045 75.510 565.275 77.390 ;
		LAYER M4 ;
		RECT 548.045 84.790 565.275 86.670 ;
		LAYER M4 ;
		RECT 548.045 45.460 565.275 47.505 ;
		LAYER M4 ;
		RECT 548.045 47.670 565.275 49.550 ;
		LAYER M4 ;
		RECT 548.045 51.135 565.275 51.275 ;
		LAYER M4 ;
		RECT 548.045 53.065 565.275 53.595 ;
		LAYER M4 ;
		RECT 548.045 253.855 565.275 253.995 ;
		LAYER M4 ;
		RECT 548.045 250.390 565.275 252.270 ;
		LAYER M4 ;
		RECT 548.045 246.505 565.275 247.035 ;
		LAYER M4 ;
		RECT 548.045 244.575 565.275 244.715 ;
		LAYER M4 ;
		RECT 548.045 248.180 565.275 250.225 ;
		LAYER M4 ;
		RECT 548.045 255.785 565.275 256.315 ;
		LAYER M4 ;
		RECT 548.045 274.345 565.275 274.875 ;
		LAYER M4 ;
		RECT 548.045 276.020 565.275 278.065 ;
		LAYER M4 ;
		RECT 548.045 278.230 565.275 280.110 ;
		LAYER M4 ;
		RECT 548.045 268.950 565.275 270.830 ;
		LAYER M4 ;
		RECT 548.045 272.415 565.275 272.555 ;
		LAYER M4 ;
		RECT 548.045 281.695 565.275 281.835 ;
		LAYER M4 ;
		RECT 548.045 263.135 565.275 263.275 ;
		LAYER M4 ;
		RECT 548.045 259.670 565.275 261.550 ;
		LAYER M4 ;
		RECT 548.045 257.460 565.275 259.505 ;
		LAYER M4 ;
		RECT 548.045 265.065 565.275 265.595 ;
		LAYER M4 ;
		RECT 548.045 266.740 565.275 268.785 ;
		LAYER M4 ;
		RECT 548.045 136.585 565.275 137.115 ;
		LAYER M4 ;
		RECT 548.045 153.215 565.275 153.355 ;
		LAYER M4 ;
		RECT 548.045 149.750 565.275 151.630 ;
		LAYER M4 ;
		RECT 548.045 147.540 565.275 149.585 ;
		LAYER M4 ;
		RECT 548.045 138.260 565.275 140.305 ;
		LAYER M4 ;
		RECT 548.045 140.470 565.275 142.350 ;
		LAYER M4 ;
		RECT 548.045 143.935 565.275 144.075 ;
		LAYER M4 ;
		RECT 548.045 145.865 565.275 146.395 ;
		LAYER M4 ;
		RECT 548.045 134.655 565.275 134.795 ;
		LAYER M4 ;
		RECT 548.045 162.495 565.275 162.635 ;
		LAYER M4 ;
		RECT 548.045 155.145 565.275 155.675 ;
		LAYER M4 ;
		RECT 548.045 159.030 565.275 160.910 ;
		LAYER M4 ;
		RECT 548.045 166.100 565.275 168.145 ;
		LAYER M4 ;
		RECT 548.045 164.425 565.275 164.955 ;
		LAYER M4 ;
		RECT 548.045 185.430 565.275 187.310 ;
		LAYER M4 ;
		RECT 548.045 198.175 565.275 198.315 ;
		LAYER M4 ;
		RECT 548.045 188.895 565.275 189.035 ;
		LAYER M1 ;
		RECT 654.555 156.335 654.735 159.695 ;
		LAYER M1 ;
		RECT 654.555 159.965 654.735 160.085 ;
		LAYER M2 ;
		RECT 654.555 160.375 654.735 160.685 ;
		LAYER M2 ;
		RECT 654.555 164.895 654.735 165.300 ;
		LAYER M4 ;
		RECT 565.275 155.145 637.535 155.640 ;
		LAYER M2 ;
		RECT 654.555 156.355 654.735 159.675 ;
		LAYER M2 ;
		RECT 654.555 167.510 654.735 168.860 ;
		LAYER M3 ;
		RECT 654.555 164.895 654.735 165.300 ;
		LAYER M4 ;
		RECT 565.275 302.185 637.535 302.680 ;
		LAYER M4 ;
		RECT 565.275 292.905 637.535 293.400 ;
		LAYER M4 ;
		RECT 565.275 283.625 637.535 284.120 ;
		LAYER M4 ;
		RECT 565.275 274.345 637.535 274.840 ;
		LAYER M4 ;
		RECT 565.275 311.465 637.535 311.960 ;
		LAYER M4 ;
		RECT 548.045 216.735 565.275 216.875 ;
		LAYER M4 ;
		RECT 548.045 156.820 565.275 158.865 ;
		LAYER M4 ;
		RECT 548.045 190.825 565.275 191.355 ;
		LAYER M4 ;
		RECT 548.045 213.270 565.275 215.150 ;
		LAYER M4 ;
		RECT 548.045 211.060 565.275 213.105 ;
		LAYER M4 ;
		RECT 548.045 192.500 565.275 194.545 ;
		LAYER M4 ;
		RECT 548.045 209.385 565.275 209.915 ;
		LAYER M4 ;
		RECT 548.045 207.455 565.275 207.595 ;
		LAYER M4 ;
		RECT 548.045 203.990 565.275 205.870 ;
		LAYER M4 ;
		RECT 548.045 194.710 565.275 196.590 ;
		LAYER M2 ;
		RECT 654.555 169.170 654.735 169.250 ;
		LAYER M4 ;
		RECT 565.275 164.425 637.535 164.920 ;
		LAYER M4 ;
		RECT 565.275 190.825 637.535 191.320 ;
		LAYER M4 ;
		RECT 565.275 200.105 637.535 200.600 ;
		LAYER M4 ;
		RECT 635.910 176.545 654.735 176.905 ;
		LAYER M4 ;
		RECT 548.045 220.340 565.275 222.385 ;
		LAYER M4 ;
		RECT 565.275 227.945 637.535 228.440 ;
		LAYER M4 ;
		RECT 565.275 237.225 637.535 237.720 ;
		LAYER M4 ;
		RECT 565.275 246.505 637.535 247.000 ;
		LAYER M4 ;
		RECT 565.275 265.065 637.535 265.560 ;
		LAYER M4 ;
		RECT 565.275 255.785 637.535 256.280 ;
		LAYER M4 ;
		RECT 565.275 218.665 637.535 219.160 ;
		LAYER M4 ;
		RECT 565.275 209.385 637.535 209.880 ;
		LAYER M4 ;
		RECT 565.275 34.505 637.535 35.000 ;
		LAYER M4 ;
		RECT 565.275 25.225 637.535 25.720 ;
		LAYER M4 ;
		RECT 565.275 15.945 637.535 16.440 ;
		LAYER M4 ;
		RECT 548.045 6.665 565.275 7.195 ;
		LAYER M4 ;
		RECT 565.275 43.785 637.535 44.280 ;
		LAYER M4 ;
		RECT 565.275 108.745 637.535 109.240 ;
		LAYER M4 ;
		RECT 548.045 108.745 565.275 109.275 ;
		LAYER M4 ;
		RECT 548.045 90.185 565.275 90.715 ;
		LAYER M4 ;
		RECT 565.275 90.185 637.535 90.680 ;
		LAYER M4 ;
		RECT 565.275 99.465 637.535 99.960 ;
		LAYER M4 ;
		RECT 565.275 62.345 637.535 62.840 ;
		LAYER M4 ;
		RECT 565.275 53.065 637.535 53.560 ;
		LAYER M4 ;
		RECT 565.275 71.625 637.535 72.120 ;
		LAYER M4 ;
		RECT 565.275 80.905 637.535 81.400 ;
		LAYER M4 ;
		RECT 548.045 62.345 565.275 62.875 ;
		LAYER M4 ;
		RECT 548.045 64.020 565.275 66.065 ;
		LAYER M4 ;
		RECT 548.045 69.695 565.275 69.835 ;
		LAYER M1 ;
		RECT 654.555 7.855 654.735 15.855 ;
		LAYER VIA3 ;
		RECT 654.555 7.875 654.735 15.835 ;
		LAYER M1 ;
		RECT 654.555 16.125 654.735 16.245 ;
		LAYER VIA3 ;
		RECT 654.555 16.535 654.735 16.845 ;
		LAYER M2 ;
		RECT 654.555 16.145 654.735 16.225 ;
		LAYER M3 ;
		RECT 654.555 16.145 654.735 16.225 ;
		LAYER M4 ;
		RECT 637.535 34.505 654.345 35.500 ;
		LAYER M4 ;
		RECT 637.535 31.670 654.345 32.715 ;
		LAYER M4 ;
		RECT 637.535 13.110 654.345 14.155 ;
		LAYER M4 ;
		RECT 637.535 15.945 654.345 16.940 ;
		LAYER M4 ;
		RECT 637.535 105.910 654.345 106.955 ;
		LAYER M4 ;
		RECT 565.275 118.025 637.535 118.520 ;
		LAYER M4 ;
		RECT 565.275 127.305 637.535 127.800 ;
		LAYER M4 ;
		RECT 565.275 136.585 637.535 137.080 ;
		LAYER M4 ;
		RECT 637.535 59.510 654.345 60.555 ;
		LAYER M4 ;
		RECT 637.535 99.465 654.345 100.460 ;
		LAYER M2 ;
		RECT 654.555 6.865 654.735 6.945 ;
		LAYER M3 ;
		RECT 654.555 6.865 654.735 6.945 ;
		LAYER VIA3 ;
		RECT 654.555 6.865 654.735 6.945 ;
		LAYER VIA3 ;
		RECT 654.555 7.255 654.735 7.565 ;
		LAYER M4 ;
		RECT 565.275 6.665 637.535 7.160 ;
		LAYER M4 ;
		RECT 637.535 6.665 654.345 7.660 ;
		LAYER M4 ;
		RECT 565.275 145.865 637.535 146.360 ;
		LAYER M1 ;
		RECT 654.555 44.975 654.735 52.975 ;
		LAYER M3 ;
		RECT 654.555 54.275 654.735 62.235 ;
		LAYER VIA3 ;
		RECT 654.555 54.275 654.735 62.235 ;
		LAYER M3 ;
		RECT 654.555 26.435 654.735 34.395 ;
		LAYER M2 ;
		RECT 654.555 44.995 654.735 52.955 ;
		LAYER M1 ;
		RECT 654.555 54.255 654.735 62.255 ;
		LAYER M1 ;
		RECT 654.555 62.525 654.735 62.645 ;
		LAYER M1 ;
		RECT 654.555 62.915 654.735 63.265 ;
		LAYER M1 ;
		RECT 654.555 53.635 654.735 53.985 ;
		LAYER M4 ;
		RECT 637.535 25.225 654.345 26.220 ;
		LAYER M1 ;
		RECT 654.555 25.405 654.735 25.525 ;
		LAYER M4 ;
		RECT 637.535 22.390 654.345 23.435 ;
		LAYER M4 ;
		RECT 637.535 71.625 654.345 72.620 ;
		LAYER M4 ;
		RECT 637.535 78.070 654.345 79.115 ;
		LAYER M4 ;
		RECT 637.535 80.905 654.345 81.900 ;
		LAYER M4 ;
		RECT 637.535 87.350 654.345 88.395 ;
		LAYER M4 ;
		RECT 637.535 62.345 654.345 63.340 ;
		LAYER M4 ;
		RECT 637.535 53.065 654.345 54.060 ;
		LAYER M4 ;
		RECT 637.535 50.230 654.345 51.275 ;
		LAYER M4 ;
		RECT 637.535 40.950 654.345 41.995 ;
		LAYER M4 ;
		RECT 637.535 43.785 654.345 44.780 ;
		LAYER M4 ;
		RECT 637.535 68.790 654.345 69.835 ;
		LAYER M4 ;
		RECT 637.535 90.185 654.345 91.180 ;
		LAYER M4 ;
		RECT 637.535 96.630 654.345 97.675 ;
		LAYER M1 ;
		RECT 654.555 238.415 654.735 246.415 ;
		LAYER M1 ;
		RECT 654.555 247.695 654.735 255.695 ;
		LAYER M1 ;
		RECT 654.555 265.635 654.735 265.985 ;
		LAYER M2 ;
		RECT 654.555 266.275 654.735 274.235 ;
		LAYER VIA3 ;
		RECT 654.555 284.215 654.735 284.525 ;
		LAYER M1 ;
		RECT 654.555 283.805 654.735 283.925 ;
		LAYER M2 ;
		RECT 654.555 275.555 654.735 283.515 ;
		LAYER VIA3 ;
		RECT 654.555 274.935 654.735 275.245 ;
		LAYER M2 ;
		RECT 654.555 283.825 654.735 283.905 ;
		LAYER M3 ;
		RECT 654.555 283.825 654.735 283.905 ;
		LAYER M2 ;
		RECT 654.555 284.835 654.735 292.795 ;
		LAYER VIA3 ;
		RECT 654.555 293.105 654.735 293.185 ;
		LAYER VIA3 ;
		RECT 654.555 274.545 654.735 274.625 ;
		LAYER M1 ;
		RECT 654.555 284.195 654.735 284.545 ;
		LAYER M4 ;
		RECT 654.345 185.890 654.735 189.035 ;
		LAYER M4 ;
		RECT 637.535 185.530 654.345 189.035 ;
		LAYER M4 ;
		RECT 637.535 190.825 654.735 193.675 ;
		LAYER M4 ;
		RECT 637.535 160.645 654.735 162.635 ;
		LAYER M4 ;
		RECT 637.535 164.425 654.735 167.275 ;
		LAYER M2 ;
		RECT 654.555 312.055 654.735 312.365 ;
		LAYER M1 ;
		RECT 654.555 312.035 654.735 312.385 ;
		LAYER M2 ;
		RECT 654.555 311.665 654.735 311.745 ;
		LAYER VIA3 ;
		RECT 654.555 311.665 654.735 311.745 ;
		LAYER M4 ;
		RECT 637.535 308.630 654.345 309.675 ;
		LAYER M4 ;
		RECT 637.535 302.185 654.345 303.180 ;
		LAYER M4 ;
		RECT 637.535 317.910 654.345 318.955 ;
		LAYER M4 ;
		RECT 637.535 311.465 654.345 312.460 ;
		LAYER M1 ;
		RECT 654.555 311.645 654.735 311.765 ;
		LAYER M3 ;
		RECT 654.555 311.665 654.735 311.745 ;
		LAYER M3 ;
		RECT 654.555 312.055 654.735 312.365 ;
		LAYER VIA3 ;
		RECT 654.555 312.055 654.735 312.365 ;
		LAYER M3 ;
		RECT 654.555 302.775 654.735 303.085 ;
		LAYER M4 ;
		RECT 637.535 252.950 654.345 253.995 ;
		LAYER M4 ;
		RECT 637.535 255.785 654.345 256.780 ;
		LAYER M4 ;
		RECT 637.535 237.225 654.345 238.220 ;
		LAYER M4 ;
		RECT 637.535 234.390 654.345 235.435 ;
		LAYER M4 ;
		RECT 637.535 243.670 654.345 244.715 ;
		LAYER M4 ;
		RECT 637.535 246.505 654.345 247.500 ;
		LAYER M4 ;
		RECT 637.535 262.230 654.345 263.275 ;
		LAYER M4 ;
		RECT 637.535 271.510 654.345 272.555 ;
		LAYER VIA3 ;
		RECT 654.555 266.275 654.735 274.235 ;
		LAYER M4 ;
		RECT 637.535 274.345 654.345 275.340 ;
		LAYER M4 ;
		RECT 637.535 299.350 654.345 300.395 ;
		LAYER M4 ;
		RECT 637.535 292.905 654.345 293.900 ;
		LAYER M4 ;
		RECT 637.535 290.070 654.345 291.115 ;
		LAYER M4 ;
		RECT 637.535 283.625 654.345 284.620 ;
		LAYER VIA3 ;
		RECT 654.555 293.495 654.735 293.805 ;
		LAYER M4 ;
		RECT 637.535 215.830 654.345 216.875 ;
		LAYER M4 ;
		RECT 637.535 209.385 654.345 210.380 ;
		LAYER M4 ;
		RECT 637.535 225.110 654.345 226.155 ;
		LAYER M4 ;
		RECT 637.535 227.945 654.345 228.940 ;
		LAYER M4 ;
		RECT 637.535 206.550 654.345 207.595 ;
		LAYER M4 ;
		RECT 637.535 218.665 654.345 219.660 ;
		LAYER M4 ;
		RECT 637.535 197.270 654.345 198.315 ;
		LAYER M4 ;
		RECT 637.535 152.310 654.345 153.355 ;
		LAYER M4 ;
		RECT 637.535 155.145 654.345 156.140 ;
		LAYER M4 ;
		RECT 637.535 133.750 654.345 134.795 ;
		LAYER M4 ;
		RECT 637.535 136.585 654.345 137.580 ;
		LAYER M4 ;
		RECT 637.535 127.305 654.345 128.300 ;
		LAYER M4 ;
		RECT 637.535 124.470 654.345 125.515 ;
		LAYER M4 ;
		RECT 637.535 200.105 654.345 201.100 ;
		LAYER M4 ;
		RECT 637.535 118.025 654.345 119.020 ;
		LAYER M4 ;
		RECT 637.535 108.745 654.345 109.740 ;
		LAYER M4 ;
		RECT 637.535 115.190 654.345 116.235 ;
		LAYER M4 ;
		RECT 637.535 145.865 654.345 146.860 ;
		LAYER M4 ;
		RECT 637.535 143.030 654.345 144.075 ;
		LAYER M1 ;
		RECT 654.555 266.255 654.735 274.255 ;
		LAYER M3 ;
		RECT 654.555 266.275 654.735 274.235 ;
		LAYER M4 ;
		RECT 637.535 265.065 654.345 266.060 ;
		LAYER M4 ;
		RECT 637.535 280.790 654.345 281.835 ;
		LAYER M4 ;
		RECT 389.275 213.270 406.505 215.150 ;
		LAYER M4 ;
		RECT 389.275 211.060 406.505 213.105 ;
		LAYER M4 ;
		RECT 389.275 235.295 406.505 235.435 ;
		LAYER M4 ;
		RECT 389.275 207.455 406.505 207.595 ;
		LAYER M4 ;
		RECT 389.275 216.735 406.505 216.875 ;
		LAYER M4 ;
		RECT 389.275 218.665 406.505 219.195 ;
		LAYER M4 ;
		RECT 389.275 227.945 406.505 228.475 ;
		LAYER M4 ;
		RECT 389.275 229.620 406.505 231.665 ;
		LAYER M4 ;
		RECT 389.275 220.340 406.505 222.385 ;
		LAYER M4 ;
		RECT 389.275 222.550 406.505 224.430 ;
		LAYER M4 ;
		RECT 389.275 190.825 406.505 191.355 ;
		LAYER M4 ;
		RECT 389.275 192.500 406.505 194.545 ;
		LAYER M4 ;
		RECT 389.275 194.710 406.505 196.590 ;
		LAYER M4 ;
		RECT 389.275 198.175 406.505 198.315 ;
		LAYER M4 ;
		RECT 389.275 201.780 406.505 203.825 ;
		LAYER M4 ;
		RECT 389.275 200.105 406.505 200.635 ;
		LAYER M4 ;
		RECT 389.275 145.865 406.505 146.395 ;
		LAYER M4 ;
		RECT 389.275 143.935 406.505 144.075 ;
		LAYER M4 ;
		RECT 389.275 320.745 406.505 321.275 ;
		LAYER M4 ;
		RECT 389.275 266.740 406.505 268.785 ;
		LAYER M4 ;
		RECT 389.275 265.065 406.505 265.595 ;
		LAYER M4 ;
		RECT 389.275 315.350 406.505 317.230 ;
		LAYER M4 ;
		RECT 389.275 285.300 406.505 287.345 ;
		LAYER M4 ;
		RECT 389.275 268.950 406.505 270.830 ;
		LAYER M4 ;
		RECT 389.275 272.415 406.505 272.555 ;
		LAYER M4 ;
		RECT 389.275 309.535 406.505 309.675 ;
		LAYER M4 ;
		RECT 389.275 303.860 406.505 305.905 ;
		LAYER M4 ;
		RECT 389.275 292.905 406.505 293.435 ;
		LAYER M4 ;
		RECT 389.275 287.510 406.505 289.390 ;
		LAYER M4 ;
		RECT 389.275 300.255 406.505 300.395 ;
		LAYER M4 ;
		RECT 389.275 296.790 406.505 298.670 ;
		LAYER M4 ;
		RECT 389.275 244.575 406.505 244.715 ;
		LAYER M4 ;
		RECT 389.275 246.505 406.505 247.035 ;
		LAYER M4 ;
		RECT 389.275 253.855 406.505 253.995 ;
		LAYER M4 ;
		RECT 389.275 257.460 406.505 259.505 ;
		LAYER M4 ;
		RECT 565.275 320.745 637.535 321.240 ;
		LAYER M4 ;
		RECT 406.505 311.465 548.045 311.960 ;
		LAYER M4 ;
		RECT 406.505 246.505 548.045 247.000 ;
		LAYER M4 ;
		RECT 548.045 320.745 565.275 321.275 ;
		LAYER M4 ;
		RECT 406.505 302.185 548.045 302.680 ;
		LAYER M4 ;
		RECT 406.505 320.745 548.045 321.240 ;
		LAYER M4 ;
		RECT 406.505 237.225 548.045 237.720 ;
		LAYER M4 ;
		RECT 406.505 227.945 548.045 228.440 ;
		LAYER M4 ;
		RECT 389.275 226.015 406.505 226.155 ;
		LAYER M4 ;
		RECT 389.275 237.225 406.505 237.755 ;
		LAYER M4 ;
		RECT 389.275 238.900 406.505 240.945 ;
		LAYER M4 ;
		RECT 247.735 227.945 389.275 228.440 ;
		LAYER M4 ;
		RECT 0.000 227.945 71.735 228.440 ;
		LAYER M4 ;
		RECT 0.000 226.485 654.345 227.565 ;
		LAYER M4 ;
		RECT 0.000 217.205 654.345 218.285 ;
		LAYER M4 ;
		RECT 406.505 218.665 548.045 219.160 ;
		LAYER M4 ;
		RECT 0.000 235.295 1.365 235.435 ;
		LAYER M4 ;
		RECT 0.000 245.045 654.345 246.125 ;
		LAYER M4 ;
		RECT 0.000 272.885 654.345 273.965 ;
		LAYER M4 ;
		RECT 0.000 282.165 654.345 283.245 ;
		LAYER M4 ;
		RECT 0.000 254.325 654.345 255.405 ;
		LAYER M4 ;
		RECT 0.000 263.605 654.345 264.685 ;
		LAYER M4 ;
		RECT 389.275 294.580 406.505 296.625 ;
		LAYER M4 ;
		RECT 406.505 292.905 548.045 293.400 ;
		LAYER M4 ;
		RECT 406.505 283.625 548.045 284.120 ;
		LAYER M4 ;
		RECT 406.505 255.785 548.045 256.280 ;
		LAYER M4 ;
		RECT 406.505 265.065 548.045 265.560 ;
		LAYER M4 ;
		RECT 406.505 274.345 548.045 274.840 ;
		LAYER M4 ;
		RECT 0.000 226.015 1.365 226.155 ;
		LAYER M4 ;
		RECT 0.000 310.005 654.345 311.085 ;
		LAYER M4 ;
		RECT 0.000 291.445 654.345 292.525 ;
		LAYER M4 ;
		RECT 0.000 300.725 654.345 301.805 ;
		LAYER M4 ;
		RECT 0.000 319.285 654.345 320.365 ;
		LAYER M4 ;
		RECT 406.505 190.825 548.045 191.320 ;
		LAYER M4 ;
		RECT 406.505 145.865 548.045 146.360 ;
		LAYER M4 ;
		RECT 406.505 155.145 548.045 155.640 ;
		LAYER M4 ;
		RECT 406.505 99.465 548.045 99.960 ;
		LAYER M4 ;
		RECT 406.505 118.025 548.045 118.520 ;
		LAYER M4 ;
		RECT 406.505 164.425 548.045 164.920 ;
		LAYER M4 ;
		RECT 389.275 140.470 406.505 142.350 ;
		LAYER M4 ;
		RECT 389.275 164.425 406.505 164.955 ;
		LAYER M4 ;
		RECT 389.275 149.750 406.505 151.630 ;
		LAYER M4 ;
		RECT 389.275 147.540 406.505 149.585 ;
		LAYER M4 ;
		RECT 389.275 138.260 406.505 140.305 ;
		LAYER M4 ;
		RECT 389.275 136.585 406.505 137.115 ;
		LAYER M4 ;
		RECT 389.275 131.190 406.505 133.070 ;
		LAYER M4 ;
		RECT 389.275 125.375 406.505 125.515 ;
		LAYER M4 ;
		RECT 389.275 119.700 406.505 121.745 ;
		LAYER M4 ;
		RECT 389.275 118.025 406.505 118.555 ;
		LAYER M4 ;
		RECT 389.275 116.095 406.505 116.235 ;
		LAYER M4 ;
		RECT 389.275 99.465 406.505 99.995 ;
		LAYER M4 ;
		RECT 389.275 156.820 406.505 158.865 ;
		LAYER M4 ;
		RECT 389.275 155.145 406.505 155.675 ;
		LAYER M4 ;
		RECT 389.275 159.030 406.505 160.910 ;
		LAYER M4 ;
		RECT 389.275 162.495 406.505 162.635 ;
		LAYER M4 ;
		RECT 354.115 184.105 388.675 185.060 ;
		LAYER M4 ;
		RECT 283.595 184.105 318.155 185.060 ;
		LAYER M4 ;
		RECT 248.875 184.105 282.895 185.060 ;
		LAYER M4 ;
		RECT 318.855 183.525 388.675 184.105 ;
		LAYER M4 ;
		RECT 318.855 184.105 353.415 185.060 ;
		LAYER M4 ;
		RECT 318.155 183.525 318.855 185.060 ;
		LAYER M4 ;
		RECT 71.135 183.525 89.565 185.060 ;
		LAYER M4 ;
		RECT 248.335 183.525 318.155 184.105 ;
		LAYER M4 ;
		RECT 230.505 185.430 247.735 187.310 ;
		LAYER M4 ;
		RECT 229.905 183.525 248.335 185.060 ;
		LAYER M4 ;
		RECT 71.735 185.430 88.965 187.310 ;
		LAYER M4 ;
		RECT 1.315 183.525 71.135 184.105 ;
		LAYER M4 ;
		RECT 389.275 188.895 406.505 189.035 ;
		LAYER M4 ;
		RECT 230.505 188.895 247.735 189.035 ;
		LAYER M4 ;
		RECT 247.735 190.825 389.275 191.320 ;
		LAYER M4 ;
		RECT 230.505 190.825 247.735 191.355 ;
		LAYER M4 ;
		RECT 71.735 194.710 88.965 196.590 ;
		LAYER M4 ;
		RECT 230.505 192.500 247.735 194.545 ;
		LAYER M4 ;
		RECT 88.965 190.825 230.505 191.320 ;
		LAYER M4 ;
		RECT 230.505 194.710 247.735 196.590 ;
		LAYER M4 ;
		RECT 389.275 153.215 406.505 153.355 ;
		LAYER M4 ;
		RECT 389.275 134.655 406.505 134.795 ;
		LAYER M4 ;
		RECT 247.735 136.585 389.275 137.080 ;
		LAYER M4 ;
		RECT 247.735 127.305 389.275 127.800 ;
		LAYER M4 ;
		RECT 247.735 155.145 389.275 155.640 ;
		LAYER M4 ;
		RECT 230.505 156.820 247.735 158.865 ;
		LAYER M4 ;
		RECT 230.505 159.030 247.735 160.910 ;
		LAYER M4 ;
		RECT 230.505 162.495 247.735 162.635 ;
		LAYER M4 ;
		RECT 230.505 155.145 247.735 155.675 ;
		LAYER M4 ;
		RECT 247.735 145.865 389.275 146.360 ;
		LAYER M4 ;
		RECT 230.505 147.540 247.735 149.585 ;
		LAYER M4 ;
		RECT 230.505 149.750 247.735 151.630 ;
		LAYER M4 ;
		RECT 71.735 166.100 88.965 168.145 ;
		LAYER M4 ;
		RECT 230.505 166.100 247.735 168.145 ;
		LAYER M4 ;
		RECT 230.505 164.425 247.735 164.955 ;
		LAYER M4 ;
		RECT 247.735 164.425 389.275 164.920 ;
		LAYER M4 ;
		RECT 88.965 108.745 230.505 109.240 ;
		LAYER M4 ;
		RECT 247.735 108.745 389.275 109.240 ;
		LAYER M4 ;
		RECT 247.735 99.465 389.275 99.960 ;
		LAYER M4 ;
		RECT 230.505 207.455 247.735 207.595 ;
		LAYER M4 ;
		RECT 230.505 203.990 247.735 205.870 ;
		LAYER M4 ;
		RECT 230.505 201.780 247.735 203.825 ;
		LAYER M4 ;
		RECT 230.505 200.105 247.735 200.635 ;
		LAYER M4 ;
		RECT 406.505 200.105 548.045 200.600 ;
		LAYER M4 ;
		RECT 230.505 198.175 247.735 198.315 ;
		LAYER M4 ;
		RECT 247.735 200.105 389.275 200.600 ;
		LAYER M4 ;
		RECT 88.965 200.105 230.505 200.600 ;
		LAYER M4 ;
		RECT 0.000 198.645 654.345 199.725 ;
		LAYER M4 ;
		RECT 0.000 209.385 71.735 209.880 ;
		LAYER M4 ;
		RECT 71.735 209.385 88.965 209.915 ;
		LAYER M4 ;
		RECT 88.965 209.385 230.505 209.880 ;
		LAYER M4 ;
		RECT 230.505 209.385 247.735 209.915 ;
		LAYER M4 ;
		RECT 406.505 209.385 548.045 209.880 ;
		LAYER M4 ;
		RECT 389.275 209.385 406.505 209.915 ;
		LAYER M4 ;
		RECT 247.735 209.385 389.275 209.880 ;
		LAYER M4 ;
		RECT 389.275 203.990 406.505 205.870 ;
		LAYER M4 ;
		RECT 0.000 207.455 1.365 207.595 ;
		LAYER M4 ;
		RECT 71.735 207.455 88.965 207.595 ;
		LAYER M4 ;
		RECT 0.000 207.925 654.345 209.005 ;
		LAYER M4 ;
		RECT 71.735 200.105 88.965 200.635 ;
		LAYER M4 ;
		RECT 71.735 198.175 88.965 198.315 ;
		LAYER M4 ;
		RECT 71.735 201.780 88.965 203.825 ;
		LAYER M4 ;
		RECT 71.735 203.990 88.965 205.870 ;
		LAYER M4 ;
		RECT 0.000 198.175 1.365 198.315 ;
		LAYER M4 ;
		RECT 71.735 108.745 88.965 109.275 ;
		LAYER M4 ;
		RECT 71.735 106.815 88.965 106.955 ;
		LAYER M4 ;
		RECT 71.735 110.420 88.965 112.465 ;
		LAYER M4 ;
		RECT 71.735 121.910 88.965 123.790 ;
		LAYER M4 ;
		RECT 0.000 108.745 71.735 109.240 ;
		LAYER M4 ;
		RECT 406.505 127.305 548.045 127.800 ;
		LAYER M4 ;
		RECT 0.000 116.565 654.345 117.645 ;
		LAYER M4 ;
		RECT 247.735 118.025 389.275 118.520 ;
		LAYER M4 ;
		RECT 0.000 107.285 654.345 108.365 ;
		LAYER M4 ;
		RECT 230.505 125.375 247.735 125.515 ;
		LAYER M4 ;
		RECT 71.735 125.375 88.965 125.515 ;
		LAYER M4 ;
		RECT 0.000 125.845 654.345 126.925 ;
		LAYER M4 ;
		RECT 71.735 155.145 88.965 155.675 ;
		LAYER M4 ;
		RECT 0.000 153.685 654.345 154.765 ;
		LAYER M4 ;
		RECT 0.000 144.405 654.345 145.485 ;
		LAYER M4 ;
		RECT 0.000 127.305 71.735 127.800 ;
		LAYER M4 ;
		RECT 71.735 127.305 88.965 127.835 ;
		LAYER M4 ;
		RECT 0.000 136.585 71.735 137.080 ;
		LAYER M4 ;
		RECT 0.000 135.125 654.345 136.205 ;
		LAYER M4 ;
		RECT 389.275 248.180 406.505 250.225 ;
		LAYER M4 ;
		RECT 389.275 311.465 406.505 311.995 ;
		LAYER M4 ;
		RECT 389.275 306.070 406.505 307.950 ;
		LAYER M4 ;
		RECT 389.275 318.815 406.505 318.955 ;
		LAYER M4 ;
		RECT 389.275 313.140 406.505 315.185 ;
		LAYER M4 ;
		RECT 389.275 250.390 406.505 252.270 ;
		LAYER M4 ;
		RECT 389.275 302.185 406.505 302.715 ;
		LAYER M4 ;
		RECT 389.275 290.975 406.505 291.115 ;
		LAYER M4 ;
		RECT 389.275 255.785 406.505 256.315 ;
		LAYER M4 ;
		RECT 389.275 259.670 406.505 261.550 ;
		LAYER M4 ;
		RECT 389.275 263.135 406.505 263.275 ;
		LAYER M4 ;
		RECT 389.275 281.695 406.505 281.835 ;
		LAYER M4 ;
		RECT 389.275 283.625 406.505 284.155 ;
		LAYER M4 ;
		RECT 230.505 296.790 247.735 298.670 ;
		LAYER M4 ;
		RECT 230.505 294.580 247.735 296.625 ;
		LAYER M4 ;
		RECT 230.505 302.185 247.735 302.715 ;
		LAYER M4 ;
		RECT 230.505 303.860 247.735 305.905 ;
		LAYER M4 ;
		RECT 230.505 300.255 247.735 300.395 ;
		LAYER M4 ;
		RECT 230.505 306.070 247.735 307.950 ;
		LAYER M4 ;
		RECT 230.505 292.905 247.735 293.435 ;
		LAYER M4 ;
		RECT 230.505 290.975 247.735 291.115 ;
		LAYER M4 ;
		RECT 230.505 287.510 247.735 289.390 ;
		LAYER M4 ;
		RECT 230.505 276.020 247.735 278.065 ;
		LAYER M4 ;
		RECT 230.505 274.345 247.735 274.875 ;
		LAYER M4 ;
		RECT 230.505 272.415 247.735 272.555 ;
		LAYER M4 ;
		RECT 230.505 266.740 247.735 268.785 ;
		LAYER M4 ;
		RECT 230.505 268.950 247.735 270.830 ;
		LAYER M4 ;
		RECT 230.505 320.745 247.735 321.275 ;
		LAYER M4 ;
		RECT 230.505 313.140 247.735 315.185 ;
		LAYER M4 ;
		RECT 230.505 265.065 247.735 265.595 ;
		LAYER M4 ;
		RECT 230.505 318.815 247.735 318.955 ;
		LAYER M4 ;
		RECT 230.505 315.350 247.735 317.230 ;
		LAYER M4 ;
		RECT 230.505 311.465 247.735 311.995 ;
		LAYER M4 ;
		RECT 230.505 278.230 247.735 280.110 ;
		LAYER M4 ;
		RECT 230.505 281.695 247.735 281.835 ;
		LAYER M4 ;
		RECT 230.505 309.535 247.735 309.675 ;
		LAYER M4 ;
		RECT 230.505 283.625 247.735 284.155 ;
		LAYER M4 ;
		RECT 230.505 285.300 247.735 287.345 ;
		LAYER M4 ;
		RECT 88.965 274.345 230.505 274.840 ;
		LAYER M4 ;
		RECT 230.505 250.390 247.735 252.270 ;
		LAYER M4 ;
		RECT 230.505 255.785 247.735 256.315 ;
		LAYER M4 ;
		RECT 88.965 265.065 230.505 265.560 ;
		LAYER M4 ;
		RECT 247.735 274.345 389.275 274.840 ;
		LAYER M4 ;
		RECT 247.735 265.065 389.275 265.560 ;
		LAYER M4 ;
		RECT 230.505 263.135 247.735 263.275 ;
		LAYER M4 ;
		RECT 230.505 257.460 247.735 259.505 ;
		LAYER M4 ;
		RECT 230.505 259.670 247.735 261.550 ;
		LAYER M4 ;
		RECT 389.275 276.020 406.505 278.065 ;
		LAYER M4 ;
		RECT 389.275 274.345 406.505 274.875 ;
		LAYER M4 ;
		RECT 389.275 278.230 406.505 280.110 ;
		LAYER M4 ;
		RECT 247.735 283.625 389.275 284.120 ;
		LAYER M4 ;
		RECT 247.735 292.905 389.275 293.400 ;
		LAYER M4 ;
		RECT 88.965 292.905 230.505 293.400 ;
		LAYER M4 ;
		RECT 247.735 311.465 389.275 311.960 ;
		LAYER M4 ;
		RECT 247.735 320.745 389.275 321.240 ;
		LAYER M4 ;
		RECT 88.965 302.185 230.505 302.680 ;
		LAYER M4 ;
		RECT 88.965 311.465 230.505 311.960 ;
		LAYER M4 ;
		RECT 88.965 320.745 230.505 321.240 ;
		LAYER M4 ;
		RECT 88.965 283.625 230.505 284.120 ;
		LAYER M4 ;
		RECT 389.275 241.110 406.505 242.990 ;
		LAYER M4 ;
		RECT 247.735 237.225 389.275 237.720 ;
		LAYER M4 ;
		RECT 247.735 246.505 389.275 247.000 ;
		LAYER M4 ;
		RECT 230.505 246.505 247.735 247.035 ;
		LAYER M4 ;
		RECT 0.000 244.575 1.365 244.715 ;
		LAYER M4 ;
		RECT 0.000 253.855 1.365 253.995 ;
		LAYER M4 ;
		RECT 0.000 246.505 71.735 247.000 ;
		LAYER M4 ;
		RECT 0.000 255.785 71.735 256.280 ;
		LAYER M4 ;
		RECT 88.965 218.665 230.505 219.160 ;
		LAYER M4 ;
		RECT 88.965 246.505 230.505 247.000 ;
		LAYER M4 ;
		RECT 88.965 237.225 230.505 237.720 ;
		LAYER M4 ;
		RECT 88.965 227.945 230.505 228.440 ;
		LAYER M4 ;
		RECT 88.965 255.785 230.505 256.280 ;
		LAYER M4 ;
		RECT 247.735 255.785 389.275 256.280 ;
		LAYER M4 ;
		RECT 247.735 218.665 389.275 219.160 ;
		LAYER M4 ;
		RECT 230.505 226.015 247.735 226.155 ;
		LAYER M4 ;
		RECT 230.505 253.855 247.735 253.995 ;
		LAYER M4 ;
		RECT 0.000 300.255 1.365 300.395 ;
		LAYER M4 ;
		RECT 0.000 309.535 1.365 309.675 ;
		LAYER M4 ;
		RECT 0.000 216.735 1.365 216.875 ;
		LAYER M4 ;
		RECT 71.735 320.745 88.965 321.275 ;
		LAYER M4 ;
		RECT 71.735 309.535 88.965 309.675 ;
		LAYER M4 ;
		RECT 71.735 268.950 88.965 270.830 ;
		LAYER M4 ;
		RECT 71.735 266.740 88.965 268.785 ;
		LAYER M4 ;
		RECT 0.000 318.815 1.365 318.955 ;
		LAYER M4 ;
		RECT 71.735 313.140 88.965 315.185 ;
		LAYER M4 ;
		RECT 0.000 311.465 71.735 311.960 ;
		LAYER M4 ;
		RECT 71.735 311.465 88.965 311.995 ;
		LAYER M4 ;
		RECT 71.735 318.815 88.965 318.955 ;
		LAYER M4 ;
		RECT 71.735 315.350 88.965 317.230 ;
		LAYER M4 ;
		RECT 0.000 320.745 71.735 321.240 ;
		LAYER M4 ;
		RECT 0.000 302.185 71.735 302.680 ;
		LAYER M4 ;
		RECT 0.000 292.905 71.735 293.400 ;
		LAYER M4 ;
		RECT 0.000 283.625 71.735 284.120 ;
		LAYER M4 ;
		RECT 0.000 265.065 71.735 265.560 ;
		LAYER M4 ;
		RECT 0.000 274.345 71.735 274.840 ;
		LAYER M4 ;
		RECT 0.000 290.975 1.365 291.115 ;
		LAYER M4 ;
		RECT 0.000 281.695 1.365 281.835 ;
		LAYER M4 ;
		RECT 0.000 272.415 1.365 272.555 ;
		LAYER M4 ;
		RECT 0.000 263.135 1.365 263.275 ;
		LAYER M4 ;
		RECT 0.000 218.665 71.735 219.160 ;
		LAYER M4 ;
		RECT 71.735 222.550 88.965 224.430 ;
		LAYER M4 ;
		RECT 71.735 229.620 88.965 231.665 ;
		LAYER M4 ;
		RECT 0.000 237.225 71.735 237.720 ;
		LAYER M4 ;
		RECT 637.535 348.585 654.345 349.580 ;
		LAYER M4 ;
		RECT 637.535 345.750 654.345 346.795 ;
		LAYER M4 ;
		RECT 637.535 339.305 654.345 340.300 ;
		LAYER M4 ;
		RECT 565.275 339.305 637.535 339.800 ;
		LAYER M4 ;
		RECT 565.275 348.585 637.535 349.080 ;
		LAYER M4 ;
		RECT 637.535 336.470 654.345 337.515 ;
		LAYER M4 ;
		RECT 548.045 346.655 565.275 346.795 ;
		LAYER M4 ;
		RECT 548.045 343.190 565.275 345.070 ;
		LAYER M4 ;
		RECT 548.045 340.980 565.275 343.025 ;
		LAYER M4 ;
		RECT 548.045 330.025 565.275 330.555 ;
		LAYER M4 ;
		RECT 565.275 330.025 637.535 330.520 ;
		LAYER M4 ;
		RECT 548.045 331.700 565.275 333.745 ;
		LAYER M4 ;
		RECT 548.045 324.630 565.275 326.510 ;
		LAYER M4 ;
		RECT 548.045 328.095 565.275 328.235 ;
		LAYER M4 ;
		RECT 637.535 327.190 654.345 328.235 ;
		LAYER M4 ;
		RECT 637.535 330.025 654.345 331.020 ;
		LAYER M4 ;
		RECT 548.045 322.420 565.275 324.465 ;
		LAYER M4 ;
		RECT 0.000 328.095 1.365 328.235 ;
		LAYER M4 ;
		RECT 0.000 337.375 1.365 337.515 ;
		LAYER M4 ;
		RECT 0.000 330.025 71.735 330.520 ;
		LAYER M4 ;
		RECT 0.000 339.305 71.735 339.800 ;
		LAYER M4 ;
		RECT 71.735 331.700 88.965 333.745 ;
		LAYER M4 ;
		RECT 71.735 339.305 88.965 339.835 ;
		LAYER M4 ;
		RECT 71.735 340.980 88.965 343.025 ;
		LAYER M4 ;
		RECT 71.735 343.190 88.965 345.070 ;
		LAYER M4 ;
		RECT 230.505 350.260 247.735 352.305 ;
		LAYER M4 ;
		RECT 71.735 350.260 88.965 352.305 ;
		LAYER M4 ;
		RECT 88.965 339.305 230.505 339.800 ;
		LAYER M4 ;
		RECT 230.505 343.190 247.735 345.070 ;
		LAYER M4 ;
		RECT 230.505 346.655 247.735 346.795 ;
		LAYER M4 ;
		RECT 88.965 330.025 230.505 330.520 ;
		LAYER M4 ;
		RECT 247.735 339.305 389.275 339.800 ;
		LAYER M4 ;
		RECT 230.505 339.305 247.735 339.835 ;
		LAYER M4 ;
		RECT 247.735 348.585 389.275 349.080 ;
		LAYER M4 ;
		RECT 230.505 340.980 247.735 343.025 ;
		LAYER M4 ;
		RECT 71.735 324.630 88.965 326.510 ;
		LAYER M4 ;
		RECT 71.735 328.095 88.965 328.235 ;
		LAYER M4 ;
		RECT 71.735 346.655 88.965 346.795 ;
		LAYER M4 ;
		RECT 230.505 333.910 247.735 335.790 ;
		LAYER M4 ;
		RECT 230.505 337.375 247.735 337.515 ;
		LAYER M4 ;
		RECT 230.505 330.025 247.735 330.555 ;
		LAYER M4 ;
		RECT 230.505 328.095 247.735 328.235 ;
		LAYER M4 ;
		RECT 247.735 330.025 389.275 330.520 ;
		LAYER M4 ;
		RECT 230.505 324.630 247.735 326.510 ;
		LAYER M4 ;
		RECT 389.275 166.100 406.505 168.145 ;
		LAYER M4 ;
		RECT 389.275 128.980 406.505 131.025 ;
		LAYER M4 ;
		RECT 389.275 127.305 406.505 127.835 ;
		LAYER M4 ;
		RECT 389.275 121.910 406.505 123.790 ;
		LAYER M4 ;
		RECT 389.275 348.585 406.505 349.115 ;
		LAYER M4 ;
		RECT 548.045 348.585 565.275 349.115 ;
		LAYER M4 ;
		RECT 548.045 350.260 565.275 352.305 ;
		LAYER M4 ;
		RECT 389.275 350.260 406.505 352.305 ;
		LAYER M4 ;
		RECT 389.275 328.095 406.505 328.235 ;
		LAYER M4 ;
		RECT 548.045 333.910 565.275 335.790 ;
		LAYER M4 ;
		RECT 548.045 337.375 565.275 337.515 ;
		LAYER M4 ;
		RECT 406.505 136.585 548.045 137.080 ;
		LAYER M4 ;
		RECT 389.275 110.420 406.505 112.465 ;
		LAYER M4 ;
		RECT 389.275 108.745 406.505 109.275 ;
		LAYER M4 ;
		RECT 389.275 106.815 406.505 106.955 ;
		LAYER M4 ;
		RECT 406.505 90.185 548.045 90.680 ;
		LAYER M4 ;
		RECT 406.505 108.745 548.045 109.240 ;
		LAYER M4 ;
		RECT 406.505 71.625 548.045 72.120 ;
		LAYER M4 ;
		RECT 406.505 80.905 548.045 81.400 ;
		LAYER M4 ;
		RECT 0.000 88.725 654.345 89.805 ;
		LAYER M4 ;
		RECT 637.535 320.745 654.345 321.740 ;
		LAYER M4 ;
		RECT 247.735 302.185 389.275 302.680 ;
		LAYER M4 ;
		RECT 389.275 231.830 406.505 233.710 ;
		LAYER M4 ;
		RECT 0.000 235.765 654.345 236.845 ;
		LAYER M4 ;
		RECT 389.275 54.740 406.505 56.785 ;
		LAYER M4 ;
		RECT 389.275 60.415 406.505 60.555 ;
		LAYER M4 ;
		RECT 389.275 62.345 406.505 62.875 ;
		LAYER M4 ;
		RECT 389.275 64.020 406.505 66.065 ;
		LAYER M4 ;
		RECT 71.735 322.420 88.965 324.465 ;
		LAYER M4 ;
		RECT 230.505 322.420 247.735 324.465 ;
		LAYER M4 ;
		RECT 0.000 328.565 654.345 329.645 ;
		LAYER M4 ;
		RECT 389.275 346.655 406.505 346.795 ;
		LAYER M4 ;
		RECT 389.275 340.980 406.505 343.025 ;
		LAYER M4 ;
		RECT 389.275 337.375 406.505 337.515 ;
		LAYER M4 ;
		RECT 389.275 333.910 406.505 335.790 ;
		LAYER M4 ;
		RECT 389.275 343.190 406.505 345.070 ;
		LAYER M4 ;
		RECT 406.505 339.305 548.045 339.800 ;
		LAYER M4 ;
		RECT 389.275 339.305 406.505 339.835 ;
		LAYER M4 ;
		RECT 389.275 331.700 406.505 333.745 ;
		LAYER M4 ;
		RECT 389.275 322.420 406.505 324.465 ;
		LAYER M4 ;
		RECT 389.275 324.630 406.505 326.510 ;
		LAYER M4 ;
		RECT 389.275 330.025 406.505 330.555 ;
		LAYER M4 ;
		RECT 406.505 330.025 548.045 330.520 ;
		LAYER M4 ;
		RECT 71.735 306.070 88.965 307.950 ;
		LAYER M4 ;
		RECT 71.735 218.665 88.965 219.195 ;
		LAYER M4 ;
		RECT 71.735 220.340 88.965 222.385 ;
		LAYER M4 ;
		RECT 71.735 303.860 88.965 305.905 ;
		LAYER M4 ;
		RECT 71.735 244.575 88.965 244.715 ;
		LAYER M4 ;
		RECT 71.735 241.110 88.965 242.990 ;
		LAYER M4 ;
		RECT 71.735 237.225 88.965 237.755 ;
		LAYER M4 ;
		RECT 71.735 235.295 88.965 235.435 ;
		LAYER M4 ;
		RECT 71.735 238.900 88.965 240.945 ;
		LAYER M4 ;
		RECT 71.735 246.505 88.965 247.035 ;
		LAYER M4 ;
		RECT 71.735 248.180 88.965 250.225 ;
		LAYER M4 ;
		RECT 71.735 250.390 88.965 252.270 ;
		LAYER M4 ;
		RECT 71.735 253.855 88.965 253.995 ;
		LAYER M4 ;
		RECT 71.735 302.185 88.965 302.715 ;
		LAYER M4 ;
		RECT 71.735 227.945 88.965 228.475 ;
		LAYER M4 ;
		RECT 71.735 226.015 88.965 226.155 ;
		LAYER M4 ;
		RECT 71.735 231.830 88.965 233.710 ;
		LAYER M4 ;
		RECT 71.735 300.255 88.965 300.395 ;
		LAYER M4 ;
		RECT 71.735 265.065 88.965 265.595 ;
		LAYER M4 ;
		RECT 71.735 278.230 88.965 280.110 ;
		LAYER M4 ;
		RECT 71.735 287.510 88.965 289.390 ;
		LAYER M4 ;
		RECT 71.735 285.300 88.965 287.345 ;
		LAYER M4 ;
		RECT 71.735 283.625 88.965 284.155 ;
		LAYER M4 ;
		RECT 71.735 281.695 88.965 281.835 ;
		LAYER M4 ;
		RECT 71.735 296.790 88.965 298.670 ;
		LAYER M4 ;
		RECT 71.735 255.785 88.965 256.315 ;
		LAYER M4 ;
		RECT 71.735 263.135 88.965 263.275 ;
		LAYER M4 ;
		RECT 71.735 257.460 88.965 259.505 ;
		LAYER M4 ;
		RECT 71.735 259.670 88.965 261.550 ;
		LAYER M4 ;
		RECT 71.735 294.580 88.965 296.625 ;
		LAYER M4 ;
		RECT 71.735 292.905 88.965 293.435 ;
		LAYER M4 ;
		RECT 71.735 290.975 88.965 291.115 ;
		LAYER M4 ;
		RECT 71.735 272.415 88.965 272.555 ;
		LAYER M4 ;
		RECT 71.735 274.345 88.965 274.875 ;
		LAYER M4 ;
		RECT 71.735 276.020 88.965 278.065 ;
		LAYER M4 ;
		RECT 71.735 118.025 88.965 118.555 ;
		LAYER M4 ;
		RECT 71.735 216.735 88.965 216.875 ;
		LAYER M4 ;
		RECT 71.735 54.740 88.965 56.785 ;
		LAYER M4 ;
		RECT 71.735 82.580 88.965 84.625 ;
		LAYER M4 ;
		RECT 71.735 88.255 88.965 88.395 ;
		LAYER M4 ;
		RECT 71.735 97.535 88.965 97.675 ;
		LAYER M4 ;
		RECT 71.735 119.700 88.965 121.745 ;
		LAYER M4 ;
		RECT 71.735 159.030 88.965 160.910 ;
		LAYER M4 ;
		RECT 71.735 211.060 88.965 213.105 ;
		LAYER M4 ;
		RECT 71.735 213.270 88.965 215.150 ;
		LAYER M4 ;
		RECT 389.275 51.135 406.505 51.275 ;
		LAYER M4 ;
		RECT 230.505 51.135 247.735 51.275 ;
		LAYER M4 ;
		RECT 389.275 91.860 406.505 93.905 ;
		LAYER M4 ;
		RECT 389.275 94.070 406.505 95.950 ;
		LAYER M4 ;
		RECT 230.505 238.900 247.735 240.945 ;
		LAYER M4 ;
		RECT 230.505 231.830 247.735 233.710 ;
		LAYER M4 ;
		RECT 230.505 229.620 247.735 231.665 ;
		LAYER M4 ;
		RECT 230.505 227.945 247.735 228.475 ;
		LAYER M4 ;
		RECT 230.505 237.225 247.735 237.755 ;
		LAYER M4 ;
		RECT 230.505 235.295 247.735 235.435 ;
		LAYER M4 ;
		RECT 230.505 241.110 247.735 242.990 ;
		LAYER M4 ;
		RECT 230.505 244.575 247.735 244.715 ;
		LAYER M4 ;
		RECT 230.505 248.180 247.735 250.225 ;
		LAYER M4 ;
		RECT 230.505 222.550 247.735 224.430 ;
		LAYER M4 ;
		RECT 230.505 220.340 247.735 222.385 ;
		LAYER M4 ;
		RECT 230.505 218.665 247.735 219.195 ;
		LAYER M4 ;
		RECT 230.505 216.735 247.735 216.875 ;
		LAYER M4 ;
		RECT 230.505 47.670 247.735 49.550 ;
		LAYER M4 ;
		RECT 230.505 211.060 247.735 213.105 ;
		LAYER M4 ;
		RECT 230.505 213.270 247.735 215.150 ;
		LAYER M4 ;
		RECT 0.000 183.525 1.315 185.060 ;
		LAYER M4 ;
		RECT 0.000 162.495 1.365 162.635 ;
		LAYER M4 ;
		RECT 71.735 156.820 88.965 158.865 ;
		LAYER M4 ;
		RECT 0.000 164.425 71.735 164.920 ;
		LAYER M4 ;
		RECT 71.735 164.425 88.965 164.955 ;
		LAYER M4 ;
		RECT 71.735 162.495 88.965 162.635 ;
		LAYER M4 ;
		RECT 71.735 190.825 88.965 191.355 ;
		LAYER M4 ;
		RECT 0.000 190.825 71.735 191.320 ;
		LAYER M4 ;
		RECT 0.000 200.105 71.735 200.600 ;
		LAYER M4 ;
		RECT 71.735 192.500 88.965 194.545 ;
		LAYER M4 ;
		RECT 195.345 184.105 229.905 185.060 ;
		LAYER M4 ;
		RECT 160.085 184.105 194.645 185.060 ;
		LAYER M4 ;
		RECT 124.825 184.105 159.385 185.060 ;
		LAYER M4 ;
		RECT 160.085 183.525 229.905 184.105 ;
		LAYER M4 ;
		RECT 90.105 184.105 124.125 185.060 ;
		LAYER M4 ;
		RECT 88.965 164.425 230.505 164.920 ;
		LAYER M4 ;
		RECT 159.385 183.525 160.085 185.060 ;
		LAYER M4 ;
		RECT 89.565 183.525 159.385 184.105 ;
		LAYER M4 ;
		RECT 0.000 188.895 1.365 189.035 ;
		LAYER M4 ;
		RECT 71.735 188.895 88.965 189.035 ;
		LAYER M4 ;
		RECT 1.315 184.105 35.875 185.060 ;
		LAYER M4 ;
		RECT 36.575 184.105 71.135 185.060 ;
		LAYER M4 ;
		RECT 230.505 82.580 247.735 84.625 ;
		LAYER M4 ;
		RECT 230.505 99.465 247.735 99.995 ;
		LAYER M4 ;
		RECT 230.505 101.140 247.735 103.185 ;
		LAYER M4 ;
		RECT 230.505 134.655 247.735 134.795 ;
		LAYER M4 ;
		RECT 230.505 127.305 247.735 127.835 ;
		LAYER M4 ;
		RECT 230.505 119.700 247.735 121.745 ;
		LAYER M4 ;
		RECT 230.505 118.025 247.735 118.555 ;
		LAYER M4 ;
		RECT 230.505 153.215 247.735 153.355 ;
		LAYER M4 ;
		RECT 230.505 143.935 247.735 144.075 ;
		LAYER M4 ;
		RECT 230.505 138.260 247.735 140.305 ;
		LAYER M4 ;
		RECT 230.505 136.585 247.735 137.115 ;
		LAYER M4 ;
		RECT 230.505 140.470 247.735 142.350 ;
		LAYER M4 ;
		RECT 230.505 145.865 247.735 146.395 ;
		LAYER M4 ;
		RECT 230.505 116.095 247.735 116.235 ;
		LAYER M4 ;
		RECT 230.505 112.630 247.735 114.510 ;
		LAYER M4 ;
		RECT 230.505 110.420 247.735 112.465 ;
		LAYER M4 ;
		RECT 230.505 103.350 247.735 105.230 ;
		LAYER M4 ;
		RECT 230.505 108.745 247.735 109.275 ;
		LAYER M4 ;
		RECT 230.505 106.815 247.735 106.955 ;
		LAYER M4 ;
		RECT 71.735 153.215 88.965 153.355 ;
		LAYER M4 ;
		RECT 71.735 149.750 88.965 151.630 ;
		LAYER M4 ;
		RECT 71.735 147.540 88.965 149.585 ;
		LAYER M4 ;
		RECT 71.735 145.865 88.965 146.395 ;
		LAYER M4 ;
		RECT 88.965 155.145 230.505 155.640 ;
		LAYER M4 ;
		RECT 0.000 125.375 1.365 125.515 ;
		LAYER M4 ;
		RECT 0.000 116.095 1.365 116.235 ;
		LAYER M4 ;
		RECT 71.735 116.095 88.965 116.235 ;
		LAYER M4 ;
		RECT 71.735 131.190 88.965 133.070 ;
		LAYER M4 ;
		RECT 71.735 128.980 88.965 131.025 ;
		LAYER M4 ;
		RECT 0.000 118.025 71.735 118.520 ;
		LAYER M4 ;
		RECT 71.735 99.465 88.965 99.995 ;
		LAYER M4 ;
		RECT 0.000 99.465 71.735 99.960 ;
		LAYER M4 ;
		RECT 71.735 140.470 88.965 142.350 ;
		LAYER M4 ;
		RECT 71.735 103.350 88.965 105.230 ;
		LAYER M4 ;
		RECT 71.735 101.140 88.965 103.185 ;
		LAYER M4 ;
		RECT 230.505 80.905 247.735 81.435 ;
		LAYER M4 ;
		RECT 88.965 80.905 230.505 81.400 ;
		LAYER M4 ;
		RECT 230.505 90.185 247.735 90.715 ;
		LAYER M4 ;
		RECT 71.735 91.860 88.965 93.905 ;
		LAYER M4 ;
		RECT 71.735 80.905 88.965 81.435 ;
		LAYER M4 ;
		RECT 0.000 80.905 71.735 81.400 ;
		LAYER M4 ;
		RECT 0.000 155.145 71.735 155.640 ;
		LAYER M4 ;
		RECT 71.735 143.935 88.965 144.075 ;
		LAYER M4 ;
		RECT 0.000 145.865 71.735 146.360 ;
		LAYER M4 ;
		RECT 0.000 153.215 1.365 153.355 ;
		LAYER M4 ;
		RECT 0.000 143.935 1.365 144.075 ;
		LAYER M4 ;
		RECT 0.000 106.815 1.365 106.955 ;
		LAYER M4 ;
		RECT 71.735 134.655 88.965 134.795 ;
		LAYER M4 ;
		RECT 71.735 136.585 88.965 137.115 ;
		LAYER M4 ;
		RECT 71.735 138.260 88.965 140.305 ;
		LAYER M4 ;
		RECT 71.735 112.630 88.965 114.510 ;
		LAYER M4 ;
		RECT 0.000 134.655 1.365 134.795 ;
		LAYER M4 ;
		RECT 230.505 78.975 247.735 79.115 ;
		LAYER M4 ;
		RECT 230.505 66.230 247.735 68.110 ;
		LAYER M4 ;
		RECT 230.505 54.740 247.735 56.785 ;
		LAYER M4 ;
		RECT 230.505 75.510 247.735 77.390 ;
		LAYER M4 ;
		RECT 230.505 73.300 247.735 75.345 ;
		LAYER M4 ;
		RECT 230.505 71.625 247.735 72.155 ;
		LAYER M4 ;
		RECT 230.505 69.695 247.735 69.835 ;
		LAYER M4 ;
		RECT 88.965 62.345 230.505 62.840 ;
		LAYER M4 ;
		RECT 88.965 71.625 230.505 72.120 ;
		LAYER M4 ;
		RECT 88.965 127.305 230.505 127.800 ;
		LAYER M4 ;
		RECT 230.505 128.980 247.735 131.025 ;
		LAYER M4 ;
		RECT 230.505 131.190 247.735 133.070 ;
		LAYER M4 ;
		RECT 88.965 118.025 230.505 118.520 ;
		LAYER M4 ;
		RECT 230.505 84.790 247.735 86.670 ;
		LAYER M4 ;
		RECT 230.505 121.910 247.735 123.790 ;
		LAYER M4 ;
		RECT 88.965 145.865 230.505 146.360 ;
		LAYER M4 ;
		RECT 88.965 99.465 230.505 99.960 ;
		LAYER M4 ;
		RECT 88.965 136.585 230.505 137.080 ;
		LAYER M4 ;
		RECT 71.735 29.110 88.965 30.990 ;
		LAYER M4 ;
		RECT 71.735 26.900 88.965 28.945 ;
		LAYER M4 ;
		RECT 71.735 36.180 88.965 38.225 ;
		LAYER M4 ;
		RECT 71.735 38.390 88.965 40.270 ;
		LAYER M4 ;
		RECT 71.735 34.505 88.965 35.035 ;
		LAYER M4 ;
		RECT 71.735 25.225 88.965 25.755 ;
		LAYER M4 ;
		RECT 71.735 53.065 88.965 53.595 ;
		LAYER M4 ;
		RECT 71.735 60.415 88.965 60.555 ;
		LAYER M4 ;
		RECT 71.735 43.785 88.965 44.315 ;
		LAYER M4 ;
		RECT 71.735 56.950 88.965 58.830 ;
		LAYER M4 ;
		RECT 71.735 17.620 88.965 19.665 ;
		LAYER M4 ;
		RECT 71.735 19.830 88.965 21.710 ;
		LAYER M4 ;
		RECT 71.735 62.345 88.965 62.875 ;
		LAYER M4 ;
		RECT 71.735 23.295 88.965 23.435 ;
		LAYER M4 ;
		RECT 0.000 43.785 71.735 44.280 ;
		LAYER M4 ;
		RECT 71.735 45.460 88.965 47.505 ;
		LAYER M4 ;
		RECT 71.735 47.670 88.965 49.550 ;
		LAYER M4 ;
		RECT 71.735 32.575 88.965 32.715 ;
		LAYER M4 ;
		RECT 0.000 25.225 71.735 25.720 ;
		LAYER M4 ;
		RECT 389.275 41.855 406.505 41.995 ;
		LAYER M4 ;
		RECT 389.275 47.670 406.505 49.550 ;
		LAYER M4 ;
		RECT 389.275 66.230 406.505 68.110 ;
		LAYER M4 ;
		RECT 389.275 43.785 406.505 44.315 ;
		LAYER M4 ;
		RECT 389.275 45.460 406.505 47.505 ;
		LAYER M4 ;
		RECT 71.735 41.855 88.965 41.995 ;
		LAYER M4 ;
		RECT 230.505 56.950 247.735 58.830 ;
		LAYER M4 ;
		RECT 230.505 60.415 247.735 60.555 ;
		LAYER M4 ;
		RECT 247.735 62.345 389.275 62.840 ;
		LAYER M4 ;
		RECT 71.735 66.230 88.965 68.110 ;
		LAYER M4 ;
		RECT 88.965 43.785 230.505 44.280 ;
		LAYER M4 ;
		RECT 88.965 53.065 230.505 53.560 ;
		LAYER M4 ;
		RECT 406.505 34.505 548.045 35.000 ;
		LAYER M4 ;
		RECT 247.735 34.505 389.275 35.000 ;
		LAYER M4 ;
		RECT 230.505 34.505 247.735 35.035 ;
		LAYER M4 ;
		RECT 230.505 53.065 247.735 53.595 ;
		LAYER M4 ;
		RECT 247.735 53.065 389.275 53.560 ;
		LAYER M4 ;
		RECT 247.735 43.785 389.275 44.280 ;
		LAYER M4 ;
		RECT 0.000 42.325 654.345 43.405 ;
		LAYER M4 ;
		RECT 406.505 43.785 548.045 44.280 ;
		LAYER M4 ;
		RECT 406.505 53.065 548.045 53.560 ;
		LAYER M4 ;
		RECT 230.505 91.860 247.735 93.905 ;
		LAYER M4 ;
		RECT 247.735 80.905 389.275 81.400 ;
		LAYER M4 ;
		RECT 0.000 60.885 654.345 61.965 ;
		LAYER M4 ;
		RECT 389.275 69.695 406.505 69.835 ;
		LAYER M4 ;
		RECT 406.505 62.345 548.045 62.840 ;
		LAYER M4 ;
		RECT 389.275 90.185 406.505 90.715 ;
		LAYER M4 ;
		RECT 247.735 90.185 389.275 90.680 ;
		LAYER M4 ;
		RECT 88.965 90.185 230.505 90.680 ;
		LAYER M4 ;
		RECT 230.505 88.255 247.735 88.395 ;
		LAYER M4 ;
		RECT 0.000 97.535 1.365 97.675 ;
		LAYER M4 ;
		RECT 71.735 94.070 88.965 95.950 ;
		LAYER M4 ;
		RECT 0.000 79.445 654.345 80.525 ;
		LAYER M4 ;
		RECT 230.505 94.070 247.735 95.950 ;
		LAYER M4 ;
		RECT 230.505 45.460 247.735 47.505 ;
		LAYER M4 ;
		RECT 230.505 41.855 247.735 41.995 ;
		LAYER M4 ;
		RECT 230.505 38.390 247.735 40.270 ;
		LAYER M4 ;
		RECT 230.505 36.180 247.735 38.225 ;
		LAYER M4 ;
		RECT 230.505 43.785 247.735 44.315 ;
		LAYER M4 ;
		RECT 230.505 64.020 247.735 66.065 ;
		LAYER M4 ;
		RECT 230.505 62.345 247.735 62.875 ;
		LAYER M4 ;
		RECT 230.505 32.575 247.735 32.715 ;
		LAYER M4 ;
		RECT 389.275 97.535 406.505 97.675 ;
		LAYER M4 ;
		RECT 230.505 97.535 247.735 97.675 ;
		LAYER M4 ;
		RECT 0.000 98.005 654.345 99.085 ;
		LAYER M4 ;
		RECT 0.000 14.015 1.365 14.155 ;
		LAYER M4 ;
		RECT 71.735 14.015 88.965 14.155 ;
		LAYER M4 ;
		RECT 0.000 15.945 71.735 16.440 ;
		LAYER M4 ;
		RECT 71.735 15.945 88.965 16.475 ;
		LAYER M4 ;
		RECT 0.000 14.485 654.345 15.565 ;
		LAYER M4 ;
		RECT 71.735 10.550 88.965 12.430 ;
		LAYER M4 ;
		RECT 230.505 10.550 247.735 12.430 ;
		LAYER M4 ;
		RECT 230.505 14.015 247.735 14.155 ;
		LAYER M4 ;
		RECT 230.505 15.945 247.735 16.475 ;
		LAYER M4 ;
		RECT 230.505 29.110 247.735 30.990 ;
		LAYER M4 ;
		RECT 88.965 25.225 230.505 25.720 ;
		LAYER M4 ;
		RECT 88.965 34.505 230.505 35.000 ;
		LAYER M4 ;
		RECT 88.965 15.945 230.505 16.440 ;
		LAYER M4 ;
		RECT 230.505 25.225 247.735 25.755 ;
		LAYER M4 ;
		RECT 230.505 26.900 247.735 28.945 ;
		LAYER M4 ;
		RECT 389.275 23.295 406.505 23.435 ;
		LAYER M4 ;
		RECT 247.735 25.225 389.275 25.720 ;
		LAYER M4 ;
		RECT 230.505 17.620 247.735 19.665 ;
		LAYER M4 ;
		RECT 230.505 23.295 247.735 23.435 ;
		LAYER M4 ;
		RECT 247.735 15.945 389.275 16.440 ;
		LAYER M4 ;
		RECT 230.505 19.830 247.735 21.710 ;
		LAYER M4 ;
		RECT 0.000 78.975 1.365 79.115 ;
		LAYER M4 ;
		RECT 0.000 60.415 1.365 60.555 ;
		LAYER M4 ;
		RECT 0.000 51.135 1.365 51.275 ;
		LAYER M4 ;
		RECT 0.000 69.695 1.365 69.835 ;
		LAYER M4 ;
		RECT 71.735 78.975 88.965 79.115 ;
		LAYER M4 ;
		RECT 71.735 75.510 88.965 77.390 ;
		LAYER M4 ;
		RECT 71.735 73.300 88.965 75.345 ;
		LAYER M4 ;
		RECT 0.000 71.625 71.735 72.120 ;
		LAYER M4 ;
		RECT 71.735 71.625 88.965 72.155 ;
		LAYER M4 ;
		RECT 0.000 62.345 71.735 62.840 ;
		LAYER M4 ;
		RECT 0.000 53.065 71.735 53.560 ;
		LAYER M4 ;
		RECT 71.735 69.695 88.965 69.835 ;
		LAYER M4 ;
		RECT 71.735 64.020 88.965 66.065 ;
		LAYER M4 ;
		RECT 0.000 88.255 1.365 88.395 ;
		LAYER M4 ;
		RECT 0.000 90.185 71.735 90.680 ;
		LAYER M4 ;
		RECT 71.735 90.185 88.965 90.715 ;
		LAYER M4 ;
		RECT 71.735 84.790 88.965 86.670 ;
		LAYER M4 ;
		RECT 548.045 1.270 565.275 3.150 ;
		LAYER M4 ;
		RECT 548.045 4.735 565.275 4.875 ;
		LAYER M4 ;
		RECT 406.505 15.945 548.045 16.440 ;
		LAYER M4 ;
		RECT 406.505 25.225 548.045 25.720 ;
		LAYER M4 ;
		RECT 389.275 1.270 406.505 3.150 ;
		LAYER M4 ;
		RECT 0.000 6.665 71.735 7.160 ;
		LAYER M4 ;
		RECT 230.505 6.665 247.735 7.195 ;
		LAYER M4 ;
		RECT 406.505 6.665 548.045 7.160 ;
		LAYER M4 ;
		RECT 230.505 8.340 247.735 10.385 ;
		LAYER M4 ;
		RECT 637.535 3.830 654.345 4.875 ;
		LAYER M4 ;
		RECT 230.505 4.735 247.735 4.875 ;
		LAYER M4 ;
		RECT 71.735 4.735 88.965 4.875 ;
		LAYER M4 ;
		RECT 230.505 1.270 247.735 3.150 ;
		LAYER M4 ;
		RECT 247.735 71.625 389.275 72.120 ;
		LAYER M4 ;
		RECT 389.275 71.625 406.505 72.155 ;
		LAYER M4 ;
		RECT 389.275 78.975 406.505 79.115 ;
		LAYER M4 ;
		RECT 0.000 70.165 654.345 71.245 ;
		LAYER M4 ;
		RECT 389.275 75.510 406.505 77.390 ;
		LAYER M4 ;
		RECT 389.275 185.430 406.505 187.310 ;
		LAYER M4 ;
		RECT 389.275 103.350 406.505 105.230 ;
		LAYER M4 ;
		RECT 389.275 101.140 406.505 103.185 ;
		LAYER M4 ;
		RECT 389.275 112.630 406.505 114.510 ;
		LAYER M4 ;
		RECT 548.045 339.305 565.275 339.835 ;
		LAYER M4 ;
		RECT 0.000 337.845 654.345 338.925 ;
		LAYER M4 ;
		RECT 0.000 347.125 654.345 348.205 ;
		LAYER M4 ;
		RECT 0.000 346.655 1.365 346.795 ;
		LAYER M4 ;
		RECT 0.000 348.585 71.735 349.080 ;
		LAYER M4 ;
		RECT 71.735 348.585 88.965 349.115 ;
		LAYER M4 ;
		RECT 406.505 348.585 548.045 349.080 ;
		LAYER M4 ;
		RECT 230.505 348.585 247.735 349.115 ;
		LAYER M4 ;
		RECT 88.965 348.585 230.505 349.080 ;
		LAYER M2 ;
		RECT 0.000 0.000 654.555 353.410 ;
		LAYER M1 ;
		RECT 0.000 0.000 654.555 353.410 ;
		LAYER M3 ;
		RECT 0.000 0.000 654.555 353.410 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 654.555 353.410 ;
	END
	# End of OBS

END TS1N28HPCPSVTB32768X36M16SWSO

END LIBRARY
