// Copyright (c) 2024 by JLSemi Inc.
// --------------------------------------------------------------------
//
//                     JLSemi
//                     Shanghai, China
//                     Name : Zhiling Guo
//                     Email: zlguo@jlsemi.com
//
// --------------------------------------------------------------------
// --------------------------------------------------------------------
//  Revision History:1.0
//  Date          By            Revision    Design Description
//---------------------------------------------------------------------
//  2024-05-06    zlguo         1.0         ASIC
// --------------------------------------------------------------------
// --------------------------------------------------------------------
`timescale 1ns/1ns
module ASIC
(
    output  wire    PAD1_ADC_DATA_1,
    output  wire    PAD2_ADC_DATA_2,
    output  wire    PAD3_ADC_DATA_3,
    output  wire    PAD4_ADC_DATA_4,
    output  wire    PAD5_ADC_DATA_5,
    output  wire    PAD6_ADC_DATA_6,
    output  wire    PAD7_ADC_DATA_7,
    output  wire    PAD8_ADC_DATA_8,
    output  wire    PAD9_ADC_DATA_9,
    output  wire    PAD10_ADC_DATA_10,
    output  wire    PAD11_ADC_DATA_11,
    output  wire    PAD12_ADC_DATA_12,
    output  wire    PAD13_ADC_DATA_13,
    output  wire    PAD14_ADC_DATA_14,
    output  wire    PAD15_ADC_DATA_15,
    output  wire    PAD16_ADC_DATA_16,
    output  wire    PAD17_ADC_DATA_17,
    output  wire    PAD18_ADC_DATA_18,
    output  wire    PAD19_ADC_DATA_VALID,
    input   wire    PAD20_RSTN,
    output  wire    PAD21_CLK_RD,
    input   wire    PAD22_MDC,
    inout   wire    PAD23_MDIO
);

    wire            CLK200M;
    wire            ADC_CLK500M;
    wire            ADC48_CLK500M;

    wire    [8:0]   ADC_DATA_0;
    wire    [8:0]   ADC_DATA_1;
    wire    [8:0]   ADC_DATA_2;
    wire    [8:0]   ADC_DATA_3;
    wire    [8:0]   ADC_DATA_4;
    wire    [8:0]   ADC_DATA_5;
    wire    [8:0]   ADC_DATA_6;
    wire    [8:0]   ADC_DATA_7;
    wire    [8:0]   ADC_DATA_8;
    wire    [8:0]   ADC_DATA_9;
    wire    [8:0]   ADC_DATA_10;
    wire    [8:0]   ADC_DATA_11;
    wire    [8:0]   ADC_DATA_12;
    wire    [8:0]   ADC_DATA_13;
    wire    [8:0]   ADC_DATA_14;
    wire    [8:0]   ADC_DATA_15;
    wire    [8:0]   ADC_DATA_16;
    wire    [8:0]   ADC_DATA_17;
    wire    [8:0]   ADC_DATA_18;
    wire    [8:0]   ADC_DATA_19;
    wire    [8:0]   ADC_DATA_20;
    wire    [8:0]   ADC_DATA_21;
    wire    [8:0]   ADC_DATA_22;
    wire    [8:0]   ADC_DATA_23;
    wire    [8:0]   ADC_DATA_24;
    wire    [8:0]   ADC_DATA_25;
    wire    [8:0]   ADC_DATA_26;
    wire    [8:0]   ADC_DATA_27;
    wire    [8:0]   ADC_DATA_28;
    wire    [8:0]   ADC_DATA_29;
    wire    [8:0]   ADC_DATA_30;
    wire    [8:0]   ADC_DATA_31;
    wire    [8:0]   ADC_DATA_32;
    wire    [8:0]   ADC_DATA_33;
    wire    [8:0]   ADC_DATA_34;
    wire    [8:0]   ADC_DATA_35;
    wire    [8:0]   ADC_DATA_36;
    wire    [8:0]   ADC_DATA_37;
    wire    [8:0]   ADC_DATA_38;
    wire    [8:0]   ADC_DATA_39;
    wire    [8:0]   ADC_DATA_40;
    wire    [8:0]   ADC_DATA_41;
    wire    [8:0]   ADC_DATA_42;
    wire    [8:0]   ADC_DATA_43;
    wire    [8:0]   ADC_DATA_44;
    wire    [8:0]   ADC_DATA_45;
    wire    [8:0]   ADC_DATA_46;
    wire    [8:0]   ADC_DATA_47;
    wire    [8:0]   ADC_DATA_48;
    wire    [8:0]   ADC_DATA_49;
    wire    [8:0]   ADC_DATA_50;
    wire    [8:0]   ADC_DATA_51;
    wire    [8:0]   ADC_DATA_52;
    wire    [8:0]   ADC_DATA_53;
    wire    [8:0]   ADC_DATA_54;
    wire    [8:0]   ADC_DATA_55;
    wire    [8:0]   ADC_DATA_56;
    wire    [8:0]   ADC_DATA_57;
    wire    [8:0]   ADC_DATA_58;
    wire    [8:0]   ADC_DATA_59;
    wire    [8:0]   ADC_DATA_60;
    wire    [8:0]   ADC_DATA_61;
    wire    [8:0]   ADC_DATA_62;
    wire    [8:0]   ADC_DATA_63;
    wire    [8:0]   ADC_DATA_64;
    wire    [8:0]   ADC_DATA_65;
    wire    [8:0]   ADC_DATA_66;
    wire    [8:0]   ADC_DATA_67;
    wire    [8:0]   ADC_DATA_68;
    wire    [8:0]   ADC_DATA_69;
    wire    [8:0]   ADC_DATA_70;
    wire    [8:0]   ADC_DATA_71;
    wire    [8:0]   ADC_DATA_72;
    wire    [8:0]   ADC_DATA_73;
    wire    [8:0]   ADC_DATA_74;
    wire    [8:0]   ADC_DATA_75;
    wire    [8:0]   ADC_DATA_76;
    wire    [8:0]   ADC_DATA_77;
    wire    [8:0]   ADC_DATA_78;
    wire    [8:0]   ADC_DATA_79;
    wire    [8:0]   ADC_DATA_80;
    wire    [8:0]   ADC_DATA_81;
    wire    [8:0]   ADC_DATA_82;
    wire    [8:0]   ADC_DATA_83;
    wire    [8:0]   ADC_DATA_84;
    wire    [8:0]   ADC_DATA_85;
    wire    [8:0]   ADC_DATA_86;
    wire    [8:0]   ADC_DATA_87;
    wire    [8:0]   ADC_DATA_88;
    wire    [8:0]   ADC_DATA_89;
    wire    [8:0]   ADC_DATA_90;
    wire    [8:0]   ADC_DATA_91;
    wire    [8:0]   ADC_DATA_92;
    wire    [8:0]   ADC_DATA_93;
    wire    [8:0]   ADC_DATA_94;
    wire    [8:0]   ADC_DATA_95;
    wire    [8:0]   ADC48_DATA_0;
    wire    [8:0]   ADC48_DATA_1;
    wire    [8:0]   ADC48_DATA_2;
    wire    [8:0]   ADC48_DATA_3;
    wire    [8:0]   ADC48_DATA_4;
    wire    [8:0]   ADC48_DATA_5;
    wire    [8:0]   ADC48_DATA_6;
    wire    [8:0]   ADC48_DATA_7;
    wire    [8:0]   ADC48_DATA_8;
    wire    [8:0]   ADC48_DATA_9;
    wire    [8:0]   ADC48_DATA_10;
    wire    [8:0]   ADC48_DATA_11;
    wire    [8:0]   ADC48_DATA_12;
    wire    [8:0]   ADC48_DATA_13;
    wire    [8:0]   ADC48_DATA_14;
    wire    [8:0]   ADC48_DATA_15;
    wire    [8:0]   ADC48_DATA_16;
    wire    [8:0]   ADC48_DATA_17;
    wire    [8:0]   ADC48_DATA_18;
    wire    [8:0]   ADC48_DATA_19;
    wire    [8:0]   ADC48_DATA_20;
    wire    [8:0]   ADC48_DATA_21;
    wire    [8:0]   ADC48_DATA_22;
    wire    [8:0]   ADC48_DATA_23;
    wire    [8:0]   ADC48_DATA_24;
    wire    [8:0]   ADC48_DATA_25;
    wire    [8:0]   ADC48_DATA_26;
    wire    [8:0]   ADC48_DATA_27;
    wire    [8:0]   ADC48_DATA_28;
    wire    [8:0]   ADC48_DATA_29;
    wire    [8:0]   ADC48_DATA_30;
    wire    [8:0]   ADC48_DATA_31;
    wire    [8:0]   ADC48_DATA_32;
    wire    [8:0]   ADC48_DATA_33;
    wire    [8:0]   ADC48_DATA_34;
    wire    [8:0]   ADC48_DATA_35;
    wire    [8:0]   ADC48_DATA_36;
    wire    [8:0]   ADC48_DATA_37;
    wire    [8:0]   ADC48_DATA_38;
    wire    [8:0]   ADC48_DATA_39;
    wire    [8:0]   ADC48_DATA_40;
    wire    [8:0]   ADC48_DATA_41;
    wire    [8:0]   ADC48_DATA_42;
    wire    [8:0]   ADC48_DATA_43;
    wire    [8:0]   ADC48_DATA_44;
    wire    [8:0]   ADC48_DATA_45;
    wire    [8:0]   ADC48_DATA_46;
    wire    [8:0]   ADC48_DATA_47;

    // Analog register
    wire    [14:0]  SAR_PVSENSOR_CNT;
    wire            BG25M_TEST_EN;
    wire            SAR_BUFFER_PD;
    wire            SAR_CKBUF_PD;
    wire            SAR_CLK_EN;
    wire            SAR_DELAY;
    wire            SAR_PU_LDOADC;
    wire            SAR_PU_SENSOR;
    wire            SAR_PVSENSOR_CNT_EN;
    wire            SAR_REVERSE;
    wire            SAR_RSTN;
    wire            SAR_SF_ST1_PD;
    wire            SAR_SKEWGEN_EN;
    wire            SAR_TEST_EN;
    wire            SAR_VREF_PD;
    wire    [15:0]  SAR_RESVD1;
    wire    [1:0]   SAR_CKBUF_ISEL;
    wire    [1:0]   SAR_ISEL;
    wire    [1:0]   SAR_REFSEL;
    wire    [1:0]   SAR_SF_ST1_ISEL;
    wire    [2:0]   BG25M_TEST_SEL;
    wire    [2:0]   SAR_CMSEL;
    wire    [2:0]   SAR_LDO_ADCSEL;
    wire    [2:0]   SAR_LDO_BUFFERSEL;
    wire    [2:0]   SAR_LDO_CKSEL;
    wire    [2:0]   SAR_TEST_SEL;
    wire    [5:0]   SAR_CKCALBUF_DELAY;
    wire    [5:0]   SAR_DAC0_COARSE;
    wire    [5:0]   SAR_DAC0_FINE;
    wire    [5:0]   SAR_DAC1_COARSE;
    wire    [5:0]   SAR_DAC1_FINE;
    wire    [5:0]   SAR_DAC2_COARSE;
    wire    [5:0]   SAR_DAC2_FINE;
    wire    [5:0]   SAR_DAC3_COARSE;
    wire    [5:0]   SAR_DAC3_FINE;
    wire    [5:0]   SAR_DAC4_COARSE;
    wire    [5:0]   SAR_DAC4_FINE;
    wire    [5:0]   SAR_DAC5_COARSE;
    wire    [5:0]   SAR_DAC5_FINE;
    wire    [5:0]   SAR_DAC6_COARSE;
    wire    [5:0]   SAR_DAC6_FINE;
    wire    [5:0]   SAR_DAC7_COARSE;
    wire    [5:0]   SAR_DAC7_FINE;

    DIGITAL_WRAPPER
    u_digital_top
    (
    // Analog-Digital interface
    .CLK200M                    (CLK200M                    ),
    .ADC_CLK500M                (ADC_CLK500M                ),
    .ADC48_CLK500M              (ADC48_CLK500M              ),

    .ADC_DATA_0                 (ADC_DATA_0                 ),
    .ADC_DATA_1                 (ADC_DATA_1                 ),
    .ADC_DATA_2                 (ADC_DATA_2                 ),
    .ADC_DATA_3                 (ADC_DATA_3                 ),
    .ADC_DATA_4                 (ADC_DATA_4                 ),
    .ADC_DATA_5                 (ADC_DATA_5                 ),
    .ADC_DATA_6                 (ADC_DATA_6                 ),
    .ADC_DATA_7                 (ADC_DATA_7                 ),
    .ADC_DATA_8                 (ADC_DATA_8                 ),
    .ADC_DATA_9                 (ADC_DATA_9                 ),
    .ADC_DATA_10                (ADC_DATA_10                ),
    .ADC_DATA_11                (ADC_DATA_11                ),
    .ADC_DATA_12                (ADC_DATA_12                ),
    .ADC_DATA_13                (ADC_DATA_13                ),
    .ADC_DATA_14                (ADC_DATA_14                ),
    .ADC_DATA_15                (ADC_DATA_15                ),
    .ADC_DATA_16                (ADC_DATA_16                ),
    .ADC_DATA_17                (ADC_DATA_17                ),
    .ADC_DATA_18                (ADC_DATA_18                ),
    .ADC_DATA_19                (ADC_DATA_19                ),
    .ADC_DATA_20                (ADC_DATA_20                ),
    .ADC_DATA_21                (ADC_DATA_21                ),
    .ADC_DATA_22                (ADC_DATA_22                ),
    .ADC_DATA_23                (ADC_DATA_23                ),
    .ADC_DATA_24                (ADC_DATA_24                ),
    .ADC_DATA_25                (ADC_DATA_25                ),
    .ADC_DATA_26                (ADC_DATA_26                ),
    .ADC_DATA_27                (ADC_DATA_27                ),
    .ADC_DATA_28                (ADC_DATA_28                ),
    .ADC_DATA_29                (ADC_DATA_29                ),
    .ADC_DATA_30                (ADC_DATA_30                ),
    .ADC_DATA_31                (ADC_DATA_31                ),
    .ADC_DATA_32                (ADC_DATA_32                ),
    .ADC_DATA_33                (ADC_DATA_33                ),
    .ADC_DATA_34                (ADC_DATA_34                ),
    .ADC_DATA_35                (ADC_DATA_35                ),
    .ADC_DATA_36                (ADC_DATA_36                ),
    .ADC_DATA_37                (ADC_DATA_37                ),
    .ADC_DATA_38                (ADC_DATA_38                ),
    .ADC_DATA_39                (ADC_DATA_39                ),
    .ADC_DATA_40                (ADC_DATA_40                ),
    .ADC_DATA_41                (ADC_DATA_41                ),
    .ADC_DATA_42                (ADC_DATA_42                ),
    .ADC_DATA_43                (ADC_DATA_43                ),
    .ADC_DATA_44                (ADC_DATA_44                ),
    .ADC_DATA_45                (ADC_DATA_45                ),
    .ADC_DATA_46                (ADC_DATA_46                ),
    .ADC_DATA_47                (ADC_DATA_47                ),
    .ADC_DATA_48                (ADC_DATA_48                ),
    .ADC_DATA_49                (ADC_DATA_49                ),
    .ADC_DATA_50                (ADC_DATA_50                ),
    .ADC_DATA_51                (ADC_DATA_51                ),
    .ADC_DATA_52                (ADC_DATA_52                ),
    .ADC_DATA_53                (ADC_DATA_53                ),
    .ADC_DATA_54                (ADC_DATA_54                ),
    .ADC_DATA_55                (ADC_DATA_55                ),
    .ADC_DATA_56                (ADC_DATA_56                ),
    .ADC_DATA_57                (ADC_DATA_57                ),
    .ADC_DATA_58                (ADC_DATA_58                ),
    .ADC_DATA_59                (ADC_DATA_59                ),
    .ADC_DATA_60                (ADC_DATA_60                ),
    .ADC_DATA_61                (ADC_DATA_61                ),
    .ADC_DATA_62                (ADC_DATA_62                ),
    .ADC_DATA_63                (ADC_DATA_63                ),
    .ADC_DATA_64                (ADC_DATA_64                ),
    .ADC_DATA_65                (ADC_DATA_65                ),
    .ADC_DATA_66                (ADC_DATA_66                ),
    .ADC_DATA_67                (ADC_DATA_67                ),
    .ADC_DATA_68                (ADC_DATA_68                ),
    .ADC_DATA_69                (ADC_DATA_69                ),
    .ADC_DATA_70                (ADC_DATA_70                ),
    .ADC_DATA_71                (ADC_DATA_71                ),
    .ADC_DATA_72                (ADC_DATA_72                ),
    .ADC_DATA_73                (ADC_DATA_73                ),
    .ADC_DATA_74                (ADC_DATA_74                ),
    .ADC_DATA_75                (ADC_DATA_75                ),
    .ADC_DATA_76                (ADC_DATA_76                ),
    .ADC_DATA_77                (ADC_DATA_77                ),
    .ADC_DATA_78                (ADC_DATA_78                ),
    .ADC_DATA_79                (ADC_DATA_79                ),
    .ADC_DATA_80                (ADC_DATA_80                ),
    .ADC_DATA_81                (ADC_DATA_81                ),
    .ADC_DATA_82                (ADC_DATA_82                ),
    .ADC_DATA_83                (ADC_DATA_83                ),
    .ADC_DATA_84                (ADC_DATA_84                ),
    .ADC_DATA_85                (ADC_DATA_85                ),
    .ADC_DATA_86                (ADC_DATA_86                ),
    .ADC_DATA_87                (ADC_DATA_87                ),
    .ADC_DATA_88                (ADC_DATA_88                ),
    .ADC_DATA_89                (ADC_DATA_89                ),
    .ADC_DATA_90                (ADC_DATA_90                ),
    .ADC_DATA_91                (ADC_DATA_91                ),
    .ADC_DATA_92                (ADC_DATA_92                ),
    .ADC_DATA_93                (ADC_DATA_93                ),
    .ADC_DATA_94                (ADC_DATA_94                ),
    .ADC_DATA_95                (ADC_DATA_95                ),
    .ADC48_DATA_0               (ADC48_DATA_0               ),
    .ADC48_DATA_1               (ADC48_DATA_1               ),
    .ADC48_DATA_2               (ADC48_DATA_2               ),
    .ADC48_DATA_3               (ADC48_DATA_3               ),
    .ADC48_DATA_4               (ADC48_DATA_4               ),
    .ADC48_DATA_5               (ADC48_DATA_5               ),
    .ADC48_DATA_6               (ADC48_DATA_6               ),
    .ADC48_DATA_7               (ADC48_DATA_7               ),
    .ADC48_DATA_8               (ADC48_DATA_8               ),
    .ADC48_DATA_9               (ADC48_DATA_9               ),
    .ADC48_DATA_10              (ADC48_DATA_10              ),
    .ADC48_DATA_11              (ADC48_DATA_11              ),
    .ADC48_DATA_12              (ADC48_DATA_12              ),
    .ADC48_DATA_13              (ADC48_DATA_13              ),
    .ADC48_DATA_14              (ADC48_DATA_14              ),
    .ADC48_DATA_15              (ADC48_DATA_15              ),
    .ADC48_DATA_16              (ADC48_DATA_16              ),
    .ADC48_DATA_17              (ADC48_DATA_17              ),
    .ADC48_DATA_18              (ADC48_DATA_18              ),
    .ADC48_DATA_19              (ADC48_DATA_19              ),
    .ADC48_DATA_20              (ADC48_DATA_20              ),
    .ADC48_DATA_21              (ADC48_DATA_21              ),
    .ADC48_DATA_22              (ADC48_DATA_22              ),
    .ADC48_DATA_23              (ADC48_DATA_23              ),
    .ADC48_DATA_24              (ADC48_DATA_24              ),
    .ADC48_DATA_25              (ADC48_DATA_25              ),
    .ADC48_DATA_26              (ADC48_DATA_26              ),
    .ADC48_DATA_27              (ADC48_DATA_27              ),
    .ADC48_DATA_28              (ADC48_DATA_28              ),
    .ADC48_DATA_29              (ADC48_DATA_29              ),
    .ADC48_DATA_30              (ADC48_DATA_30              ),
    .ADC48_DATA_31              (ADC48_DATA_31              ),
    .ADC48_DATA_32              (ADC48_DATA_32              ),
    .ADC48_DATA_33              (ADC48_DATA_33              ),
    .ADC48_DATA_34              (ADC48_DATA_34              ),
    .ADC48_DATA_35              (ADC48_DATA_35              ),
    .ADC48_DATA_36              (ADC48_DATA_36              ),
    .ADC48_DATA_37              (ADC48_DATA_37              ),
    .ADC48_DATA_38              (ADC48_DATA_38              ),
    .ADC48_DATA_39              (ADC48_DATA_39              ),
    .ADC48_DATA_40              (ADC48_DATA_40              ),
    .ADC48_DATA_41              (ADC48_DATA_41              ),
    .ADC48_DATA_42              (ADC48_DATA_42              ),
    .ADC48_DATA_43              (ADC48_DATA_43              ),
    .ADC48_DATA_44              (ADC48_DATA_44              ),
    .ADC48_DATA_45              (ADC48_DATA_45              ),
    .ADC48_DATA_46              (ADC48_DATA_46              ),
    .ADC48_DATA_47              (ADC48_DATA_47              ),

    // Analog register
    .SAR_PVSENSOR_CNT           (SAR_PVSENSOR_CNT           ),
    .BG25M_TEST_EN              (BG25M_TEST_EN              ),
    .SAR_BUFFER_PD              (SAR_BUFFER_PD              ),
    .SAR_CKBUF_PD               (SAR_CKBUF_PD               ),
    .SAR_CLK_EN                 (SAR_CLK_EN                 ),
    .SAR_DELAY                  (SAR_DELAY                  ),
    .SAR_PU_LDOADC              (SAR_PU_LDOADC              ),
    .SAR_PU_SENSOR              (SAR_PU_SENSOR              ),
    .SAR_PVSENSOR_CNT_EN        (SAR_PVSENSOR_CNT_EN        ),
    .SAR_REVERSE                (SAR_REVERSE                ),
    .SAR_RSTN                   (SAR_RSTN                   ),
    .SAR_SF_ST1_PD              (SAR_SF_ST1_PD              ),
    .SAR_SKEWGEN_EN             (SAR_SKEWGEN_EN             ),
    .SAR_TEST_EN                (SAR_TEST_EN                ),
    .SAR_VREF_PD                (SAR_VREF_PD                ),
    .SAR_RESVD1                 (SAR_RESVD1                 ),
    .SAR_CKBUF_ISEL             (SAR_CKBUF_ISEL             ),
    .SAR_ISEL                   (SAR_ISEL                   ),
    .SAR_REFSEL                 (SAR_REFSEL                 ),
    .SAR_SF_ST1_ISEL            (SAR_SF_ST1_ISEL            ),
    .BG25M_TEST_SEL             (BG25M_TEST_SEL             ),
    .SAR_CMSEL                  (SAR_CMSEL                  ),
    .SAR_LDO_ADCSEL             (SAR_LDO_ADCSEL             ),
    .SAR_LDO_BUFFERSEL          (SAR_LDO_BUFFERSEL          ),
    .SAR_LDO_CKSEL              (SAR_LDO_CKSEL              ),
    .SAR_TEST_SEL               (SAR_TEST_SEL               ),
    .SAR_CKCALBUF_DELAY         (SAR_CKCALBUF_DELAY         ),
    .SAR_DAC0_COARSE            (SAR_DAC0_COARSE            ),
    .SAR_DAC0_FINE              (SAR_DAC0_FINE              ),
    .SAR_DAC1_COARSE            (SAR_DAC1_COARSE            ),
    .SAR_DAC1_FINE              (SAR_DAC1_FINE              ),
    .SAR_DAC2_COARSE            (SAR_DAC2_COARSE            ),
    .SAR_DAC2_FINE              (SAR_DAC2_FINE              ),
    .SAR_DAC3_COARSE            (SAR_DAC3_COARSE            ),
    .SAR_DAC3_FINE              (SAR_DAC3_FINE              ),
    .SAR_DAC4_COARSE            (SAR_DAC4_COARSE            ),
    .SAR_DAC4_FINE              (SAR_DAC4_FINE              ),
    .SAR_DAC5_COARSE            (SAR_DAC5_COARSE            ),
    .SAR_DAC5_FINE              (SAR_DAC5_FINE              ),
    .SAR_DAC6_COARSE            (SAR_DAC6_COARSE            ),
    .SAR_DAC6_FINE              (SAR_DAC6_FINE              ),
    .SAR_DAC7_COARSE            (SAR_DAC7_COARSE            ),
    .SAR_DAC7_FINE              (SAR_DAC7_FINE              ),

    // Digital io pad
    .PAD1_ADC_DATA_1            (PAD1_ADC_DATA_1            ),
    .PAD2_ADC_DATA_2            (PAD2_ADC_DATA_2            ),
    .PAD3_ADC_DATA_3            (PAD3_ADC_DATA_3            ),
    .PAD4_ADC_DATA_4            (PAD4_ADC_DATA_4            ),
    .PAD5_ADC_DATA_5            (PAD5_ADC_DATA_5            ),
    .PAD6_ADC_DATA_6            (PAD6_ADC_DATA_6            ),
    .PAD7_ADC_DATA_7            (PAD7_ADC_DATA_7            ),
    .PAD8_ADC_DATA_8            (PAD8_ADC_DATA_8            ),
    .PAD9_ADC_DATA_9            (PAD9_ADC_DATA_9            ),
    .PAD10_ADC_DATA_10          (PAD10_ADC_DATA_10          ),
    .PAD11_ADC_DATA_11          (PAD11_ADC_DATA_11          ),
    .PAD12_ADC_DATA_12          (PAD12_ADC_DATA_12          ),
    .PAD13_ADC_DATA_13          (PAD13_ADC_DATA_13          ),
    .PAD14_ADC_DATA_14          (PAD14_ADC_DATA_14          ),
    .PAD15_ADC_DATA_15          (PAD15_ADC_DATA_15          ),
    .PAD16_ADC_DATA_16          (PAD16_ADC_DATA_16          ),
    .PAD17_ADC_DATA_17          (PAD17_ADC_DATA_17          ),
    .PAD18_ADC_DATA_18          (PAD18_ADC_DATA_18          ),
    .PAD19_ADC_DATA_VALID       (PAD19_ADC_DATA_VALID       ),
    .PAD20_RSTN                 (PAD20_RSTN                 ),
    .PAD21_CLK_RD               (PAD21_CLK_RD               ),
    .PAD22_MDC                  (PAD22_MDC                  ),
    .PAD23_MDIO                 (PAD23_MDIO                 )
    );

    ANALOG_WRAPPER
    u_analog_top
    (
    // Analog to dig clock port
    .SAR_200M_REG_CLK           (CLK200M                    ),
    .HSAR_CLK_ASSO              (ADC_CLK500M                ),
    .SAR_CLK_ASSO               (ADC48_CLK500M              ),

    // Analog adc48 port
    .HSAR_DATA_0_0              (ADC_DATA_0                 ),
    .HSAR_DATA_0_1              (ADC_DATA_1                 ),
    .HSAR_DATA_0_2              (ADC_DATA_2                 ),
    .HSAR_DATA_0_3              (ADC_DATA_3                 ),
    .HSAR_DATA_0_4              (ADC_DATA_4                 ),
    .HSAR_DATA_0_5              (ADC_DATA_5                 ),
    .HSAR_DATA_0_6              (ADC_DATA_6                 ),
    .HSAR_DATA_0_7              (ADC_DATA_7                 ),
    .HSAR_DATA_0_8              (ADC_DATA_8                 ),
    .HSAR_DATA_0_9              (ADC_DATA_9                 ),
    .HSAR_DATA_1_0              (ADC_DATA_10                ),
    .HSAR_DATA_1_1              (ADC_DATA_11                ),
    .HSAR_DATA_1_2              (ADC_DATA_12                ),
    .HSAR_DATA_1_3              (ADC_DATA_13                ),
    .HSAR_DATA_1_4              (ADC_DATA_14                ),
    .HSAR_DATA_1_5              (ADC_DATA_15                ),
    .HSAR_DATA_1_6              (ADC_DATA_16                ),
    .HSAR_DATA_1_7              (ADC_DATA_17                ),
    .HSAR_DATA_1_8              (ADC_DATA_18                ),
    .HSAR_DATA_1_9              (ADC_DATA_19                ),
    .HSAR_DATA_2_0              (ADC_DATA_20                ),
    .HSAR_DATA_2_1              (ADC_DATA_21                ),
    .HSAR_DATA_2_2              (ADC_DATA_22                ),
    .HSAR_DATA_2_3              (ADC_DATA_23                ),
    .HSAR_DATA_2_4              (ADC_DATA_24                ),
    .HSAR_DATA_2_5              (ADC_DATA_25                ),
    .HSAR_DATA_2_6              (ADC_DATA_26                ),
    .HSAR_DATA_2_7              (ADC_DATA_27                ),
    .HSAR_DATA_2_8              (ADC_DATA_28                ),
    .HSAR_DATA_2_9              (ADC_DATA_29                ),
    .HSAR_DATA_3_0              (ADC_DATA_30                ),
    .HSAR_DATA_3_1              (ADC_DATA_31                ),
    .HSAR_DATA_3_2              (ADC_DATA_32                ),
    .HSAR_DATA_3_3              (ADC_DATA_33                ),
    .HSAR_DATA_3_4              (ADC_DATA_34                ),
    .HSAR_DATA_3_5              (ADC_DATA_35                ),
    .HSAR_DATA_3_6              (ADC_DATA_36                ),
    .HSAR_DATA_3_7              (ADC_DATA_37                ),
    .HSAR_DATA_3_8              (ADC_DATA_38                ),
    .HSAR_DATA_3_9              (ADC_DATA_39                ),
    .HSAR_DATA_4_0              (ADC_DATA_40                ),
    .HSAR_DATA_4_1              (ADC_DATA_41                ),
    .HSAR_DATA_4_2              (ADC_DATA_42                ),
    .HSAR_DATA_4_3              (ADC_DATA_43                ),
    .HSAR_DATA_4_4              (ADC_DATA_44                ),
    .HSAR_DATA_4_5              (ADC_DATA_45                ),
    .HSAR_DATA_4_6              (ADC_DATA_46                ),
    .HSAR_DATA_4_7              (ADC_DATA_47                ),
    .HSAR_DATA_4_8              (ADC_DATA_48                ),
    .HSAR_DATA_4_9              (ADC_DATA_49                ),
    .HSAR_DATA_5_0              (ADC_DATA_50                ),
    .HSAR_DATA_5_1              (ADC_DATA_51                ),
    .HSAR_DATA_5_2              (ADC_DATA_52                ),
    .HSAR_DATA_5_3              (ADC_DATA_53                ),
    .HSAR_DATA_5_4              (ADC_DATA_54                ),
    .HSAR_DATA_5_5              (ADC_DATA_55                ),
    .HSAR_DATA_5_6              (ADC_DATA_56                ),
    .HSAR_DATA_5_7              (ADC_DATA_57                ),
    .HSAR_DATA_5_8              (ADC_DATA_58                ),
    .HSAR_DATA_5_9              (ADC_DATA_59                ),
    .HSAR_DATA_6_0              (ADC_DATA_60                ),
    .HSAR_DATA_6_1              (ADC_DATA_61                ),
    .HSAR_DATA_6_2              (ADC_DATA_62                ),
    .HSAR_DATA_6_3              (ADC_DATA_63                ),
    .HSAR_DATA_6_4              (ADC_DATA_64                ),
    .HSAR_DATA_6_5              (ADC_DATA_65                ),
    .HSAR_DATA_6_6              (ADC_DATA_66                ),
    .HSAR_DATA_6_7              (ADC_DATA_67                ),
    .HSAR_DATA_6_8              (ADC_DATA_68                ),
    .HSAR_DATA_6_9              (ADC_DATA_69                ),
    .HSAR_DATA_7_0              (ADC_DATA_70                ),
    .HSAR_DATA_7_1              (ADC_DATA_71                ),
    .HSAR_DATA_7_2              (ADC_DATA_72                ),
    .HSAR_DATA_7_3              (ADC_DATA_73                ),
    .HSAR_DATA_7_4              (ADC_DATA_74                ),
    .HSAR_DATA_7_5              (ADC_DATA_75                ),
    .HSAR_DATA_7_6              (ADC_DATA_76                ),
    .HSAR_DATA_7_7              (ADC_DATA_77                ),
    .HSAR_DATA_7_8              (ADC_DATA_78                ),
    .HSAR_DATA_7_9              (ADC_DATA_79                ),
    .HSAR_DATA_8_0              (ADC_DATA_80                ),
    .HSAR_DATA_8_1              (ADC_DATA_81                ),
    .HSAR_DATA_8_2              (ADC_DATA_82                ),
    .HSAR_DATA_8_3              (ADC_DATA_83                ),
    .HSAR_DATA_8_4              (ADC_DATA_84                ),
    .HSAR_DATA_8_5              (ADC_DATA_85                ),
    .HSAR_DATA_8_6              (ADC_DATA_86                ),
    .HSAR_DATA_8_7              (ADC_DATA_87                ),
    .HSAR_DATA_8_8              (ADC_DATA_88                ),
    .HSAR_DATA_8_9              (ADC_DATA_89                ),
    .HSAR_DATA_9_0              (ADC_DATA_90                ),
    .HSAR_DATA_9_1              (ADC_DATA_91                ),
    .HSAR_DATA_9_2              (ADC_DATA_92                ),
    .HSAR_DATA_9_3              (ADC_DATA_93                ),
    .HSAR_DATA_9_4              (ADC_DATA_94                ),
    .HSAR_DATA_9_5              (ADC_DATA_95                ),

    // Analog adc48 port
    .SAR_DATA_0_0               (ADC48_DATA_0               ),
    .SAR_DATA_0_1               (ADC48_DATA_1               ),
    .SAR_DATA_0_2               (ADC48_DATA_2               ),
    .SAR_DATA_0_3               (ADC48_DATA_3               ),
    .SAR_DATA_0_4               (ADC48_DATA_4               ),
    .SAR_DATA_0_5               (ADC48_DATA_5               ),
    .SAR_DATA_0_6               (ADC48_DATA_6               ),
    .SAR_DATA_0_7               (ADC48_DATA_7               ),
    .SAR_DATA_0_8               (ADC48_DATA_8               ),
    .SAR_DATA_0_9               (ADC48_DATA_9               ),
    .SAR_DATA_1_0               (ADC48_DATA_10              ),
    .SAR_DATA_1_1               (ADC48_DATA_11              ),
    .SAR_DATA_1_2               (ADC48_DATA_12              ),
    .SAR_DATA_1_3               (ADC48_DATA_13              ),
    .SAR_DATA_1_4               (ADC48_DATA_14              ),
    .SAR_DATA_1_5               (ADC48_DATA_15              ),
    .SAR_DATA_1_6               (ADC48_DATA_16              ),
    .SAR_DATA_1_7               (ADC48_DATA_17              ),
    .SAR_DATA_1_8               (ADC48_DATA_18              ),
    .SAR_DATA_1_9               (ADC48_DATA_19              ),
    .SAR_DATA_2_0               (ADC48_DATA_20              ),
    .SAR_DATA_2_1               (ADC48_DATA_21              ),
    .SAR_DATA_2_2               (ADC48_DATA_22              ),
    .SAR_DATA_2_3               (ADC48_DATA_23              ),
    .SAR_DATA_2_4               (ADC48_DATA_24              ),
    .SAR_DATA_2_5               (ADC48_DATA_25              ),
    .SAR_DATA_2_6               (ADC48_DATA_26              ),
    .SAR_DATA_2_7               (ADC48_DATA_27              ),
    .SAR_DATA_2_8               (ADC48_DATA_28              ),
    .SAR_DATA_2_9               (ADC48_DATA_29              ),
    .SAR_DATA_3_0               (ADC48_DATA_30              ),
    .SAR_DATA_3_1               (ADC48_DATA_31              ),
    .SAR_DATA_3_2               (ADC48_DATA_32              ),
    .SAR_DATA_3_3               (ADC48_DATA_33              ),
    .SAR_DATA_3_4               (ADC48_DATA_34              ),
    .SAR_DATA_3_5               (ADC48_DATA_35              ),
    .SAR_DATA_3_6               (ADC48_DATA_36              ),
    .SAR_DATA_3_7               (ADC48_DATA_37              ),
    .SAR_DATA_3_8               (ADC48_DATA_38              ),
    .SAR_DATA_3_9               (ADC48_DATA_39              ),
    .SAR_DATA_4_0               (ADC48_DATA_40              ),
    .SAR_DATA_4_1               (ADC48_DATA_41              ),
    .SAR_DATA_4_2               (ADC48_DATA_42              ),
    .SAR_DATA_4_3               (ADC48_DATA_43              ),
    .SAR_DATA_4_4               (ADC48_DATA_44              ),
    .SAR_DATA_4_5               (ADC48_DATA_45              ),
    .SAR_DATA_4_6               (ADC48_DATA_46              ),
    .SAR_DATA_4_7               (ADC48_DATA_47              ),

    // Analog adc48 register
    .SAR_PVSENSOR_CNT           (SAR_PVSENSOR_CNT           ),
    .BG25M_TEST_EN              (BG25M_TEST_EN              ),
    .SAR_BUFFER_PD              (SAR_BUFFER_PD              ),
    .SAR_CKBUF_PD               (SAR_CKBUF_PD               ),
    .SAR_CLK_EN                 (SAR_CLK_EN                 ),
    .SAR_DELAY                  (SAR_DELAY                  ),
    .SAR_PU_LDOADC              (SAR_PU_LDOADC              ),
    .SAR_PU_SENSOR              (SAR_PU_SENSOR              ),
    .SAR_PVSENSOR_CNT_EN        (SAR_PVSENSOR_CNT_EN        ),
    .SAR_REVERSE                (SAR_REVERSE                ),
    .SAR_RSTN                   (SAR_RSTN                   ),
    .SAR_SF_ST1_PD              (SAR_SF_ST1_PD              ),
    .SAR_SKEWGEN_EN             (SAR_SKEWGEN_EN             ),
    .SAR_TEST_EN                (SAR_TEST_EN                ),
    .SAR_VREF_PD                (SAR_VREF_PD                ),
    .SAR_RESVD1                 (SAR_RESVD1                 ),
    .SAR_CKBUF_ISEL             (SAR_CKBUF_ISEL             ),
    .SAR_ISEL                   (SAR_ISEL                   ),
    .SAR_REFSEL                 (SAR_REFSEL                 ),
    .SAR_SF_ST1_ISEL            (SAR_SF_ST1_ISEL            ),
    .BG25M_TEST_SEL             (BG25M_TEST_SEL             ),
    .SAR_CMSEL                  (SAR_CMSEL                  ),
    .SAR_LDO_ADCSEL             (SAR_LDO_ADCSEL             ),
    .SAR_LDO_BUFFERSEL          (SAR_LDO_BUFFERSEL          ),
    .SAR_LDO_CKSEL              (SAR_LDO_CKSEL              ),
    .SAR_TEST_SEL               (SAR_TEST_SEL               ),
    .SAR_CKCALBUF_DELAY         (SAR_CKCALBUF_DELAY         ),
    .SAR_DAC0_COARSE            (SAR_DAC0_COARSE            ),
    .SAR_DAC0_FINE              (SAR_DAC0_FINE              ),
    .SAR_DAC1_COARSE            (SAR_DAC1_COARSE            ),
    .SAR_DAC1_FINE              (SAR_DAC1_FINE              ),
    .SAR_DAC2_COARSE            (SAR_DAC2_COARSE            ),
    .SAR_DAC2_FINE              (SAR_DAC2_FINE              ),
    .SAR_DAC3_COARSE            (SAR_DAC3_COARSE            ),
    .SAR_DAC3_FINE              (SAR_DAC3_FINE              ),
    .SAR_DAC4_COARSE            (SAR_DAC4_COARSE            ),
    .SAR_DAC4_FINE              (SAR_DAC4_FINE              ),
    .SAR_DAC5_COARSE            (SAR_DAC5_COARSE            ),
    .SAR_DAC5_FINE              (SAR_DAC5_FINE              ),
    .SAR_DAC6_COARSE            (SAR_DAC6_COARSE            ),
    .SAR_DAC6_FINE              (SAR_DAC6_FINE              ),
    .SAR_DAC7_COARSE            (SAR_DAC7_COARSE            ),
    .SAR_DAC7_FINE              (SAR_DAC7_FINE              ),

    .SAR_VINP                   (SAR_VINP                   ),
    .SAR_VINN                   (SAR_VINN                   ),
    .SAR_CLK_12G_IN             (SAR_CLK_12G_IN             ),
    .SAR_CLK_200M               (SAR_CLK_200M               ),
    .SAR_DVDD09                 (SAR_DVDD09                 ),
    .SAR_AVDD25_BUF             (SAR_AVDD25_BUF             ),
    .SAR_AVDD25_CK              (SAR_AVDD25_CK              ),
    .SAR_AVDD25_ADC             (SAR_AVDD25_ADC             ),
    .SAR_AVDD25                 (SAR_AVDD25                 ),
    .SAR_AGND                   (SAR_AGND                   ),
    .SAR_DVSS                   (SAR_DVSS                   ),
    .SAR_ATEST                  (SAR_ATEST                  )

    );

endmodule
