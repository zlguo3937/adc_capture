module ANALOG_WRAPPER
(
    output  wire            CLK200M,
    output  wire            CLK500M,

    output  wire    [8:0]   ADC_DATA_0,
    output  wire    [8:0]   ADC_DATA_1,
    output  wire    [8:0]   ADC_DATA_2,
    output  wire    [8:0]   ADC_DATA_3,
    output  wire    [8:0]   ADC_DATA_4,
    output  wire    [8:0]   ADC_DATA_5,
    output  wire    [8:0]   ADC_DATA_6,
    output  wire    [8:0]   ADC_DATA_7,
    output  wire    [8:0]   ADC_DATA_8,
    output  wire    [8:0]   ADC_DATA_9,
    output  wire    [8:0]   ADC_DATA_10,
    output  wire    [8:0]   ADC_DATA_11,
    output  wire    [8:0]   ADC_DATA_12,
    output  wire    [8:0]   ADC_DATA_13,
    output  wire    [8:0]   ADC_DATA_14,
    output  wire    [8:0]   ADC_DATA_15,
    output  wire    [8:0]   ADC_DATA_16,
    output  wire    [8:0]   ADC_DATA_17,
    output  wire    [8:0]   ADC_DATA_18,
    output  wire    [8:0]   ADC_DATA_19,
    output  wire    [8:0]   ADC_DATA_20,
    output  wire    [8:0]   ADC_DATA_21,
    output  wire    [8:0]   ADC_DATA_22,
    output  wire    [8:0]   ADC_DATA_23,
    output  wire    [8:0]   ADC_DATA_24,
    output  wire    [8:0]   ADC_DATA_25,
    output  wire    [8:0]   ADC_DATA_26,
    output  wire    [8:0]   ADC_DATA_27,
    output  wire    [8:0]   ADC_DATA_28,
    output  wire    [8:0]   ADC_DATA_29,
    output  wire    [8:0]   ADC_DATA_30,
    output  wire    [8:0]   ADC_DATA_31,
    output  wire    [8:0]   ADC_DATA_32,
    output  wire    [8:0]   ADC_DATA_33,
    output  wire    [8:0]   ADC_DATA_34,
    output  wire    [8:0]   ADC_DATA_35,
    output  wire    [8:0]   ADC_DATA_36,
    output  wire    [8:0]   ADC_DATA_37,
    output  wire    [8:0]   ADC_DATA_38,
    output  wire    [8:0]   ADC_DATA_39,
    output  wire    [8:0]   ADC_DATA_40,
    output  wire    [8:0]   ADC_DATA_41,
    output  wire    [8:0]   ADC_DATA_42,
    output  wire    [8:0]   ADC_DATA_43,
    output  wire    [8:0]   ADC_DATA_44,
    output  wire    [8:0]   ADC_DATA_45,
    output  wire    [8:0]   ADC_DATA_46,
    output  wire    [8:0]   ADC_DATA_47,
    output  wire    [8:0]   ADC_DATA_48,
    output  wire    [8:0]   ADC_DATA_49,
    output  wire    [8:0]   ADC_DATA_50,
    output  wire    [8:0]   ADC_DATA_51,
    output  wire    [8:0]   ADC_DATA_52,
    output  wire    [8:0]   ADC_DATA_53,
    output  wire    [8:0]   ADC_DATA_54,
    output  wire    [8:0]   ADC_DATA_55,
    output  wire    [8:0]   ADC_DATA_56,
    output  wire    [8:0]   ADC_DATA_57,
    output  wire    [8:0]   ADC_DATA_58,
    output  wire    [8:0]   ADC_DATA_59,
    output  wire    [8:0]   ADC_DATA_60,
    output  wire    [8:0]   ADC_DATA_61,
    output  wire    [8:0]   ADC_DATA_62,
    output  wire    [8:0]   ADC_DATA_63,
    output  wire    [8:0]   ADC_DATA_64,
    output  wire    [8:0]   ADC_DATA_65,
    output  wire    [8:0]   ADC_DATA_66,
    output  wire    [8:0]   ADC_DATA_67,
    output  wire    [8:0]   ADC_DATA_68,
    output  wire    [8:0]   ADC_DATA_69,
    output  wire    [8:0]   ADC_DATA_70,
    output  wire    [8:0]   ADC_DATA_71,
    output  wire    [8:0]   ADC_DATA_72,
    output  wire    [8:0]   ADC_DATA_73,
    output  wire    [8:0]   ADC_DATA_74,
    output  wire    [8:0]   ADC_DATA_75,
    output  wire    [8:0]   ADC_DATA_76,
    output  wire    [8:0]   ADC_DATA_77,
    output  wire    [8:0]   ADC_DATA_78,
    output  wire    [8:0]   ADC_DATA_79,
    output  wire    [8:0]   ADC_DATA_80,
    output  wire    [8:0]   ADC_DATA_81,
    output  wire    [8:0]   ADC_DATA_82,
    output  wire    [8:0]   ADC_DATA_83,
    output  wire    [8:0]   ADC_DATA_84,
    output  wire    [8:0]   ADC_DATA_85,
    output  wire    [8:0]   ADC_DATA_86,
    output  wire    [8:0]   ADC_DATA_87,
    output  wire    [8:0]   ADC_DATA_88,
    output  wire    [8:0]   ADC_DATA_89,
    output  wire    [8:0]   ADC_DATA_90,
    output  wire    [8:0]   ADC_DATA_91,
    output  wire    [8:0]   ADC_DATA_92,
    output  wire    [8:0]   ADC_DATA_93,
    output  wire    [8:0]   ADC_DATA_94,
    output  wire    [8:0]   ADC_DATA_95,
    output  wire    [8:0]   ADC48_DATA_0,
    output  wire    [8:0]   ADC48_DATA_1,
    output  wire    [8:0]   ADC48_DATA_2,
    output  wire    [8:0]   ADC48_DATA_3,
    output  wire    [8:0]   ADC48_DATA_4,
    output  wire    [8:0]   ADC48_DATA_5,
    output  wire    [8:0]   ADC48_DATA_6,
    output  wire    [8:0]   ADC48_DATA_7,
    output  wire    [8:0]   ADC48_DATA_8,
    output  wire    [8:0]   ADC48_DATA_9,
    output  wire    [8:0]   ADC48_DATA_10,
    output  wire    [8:0]   ADC48_DATA_11,
    output  wire    [8:0]   ADC48_DATA_12,
    output  wire    [8:0]   ADC48_DATA_13,
    output  wire    [8:0]   ADC48_DATA_14,
    output  wire    [8:0]   ADC48_DATA_15,
    output  wire    [8:0]   ADC48_DATA_16,
    output  wire    [8:0]   ADC48_DATA_17,
    output  wire    [8:0]   ADC48_DATA_18,
    output  wire    [8:0]   ADC48_DATA_19,
    output  wire    [8:0]   ADC48_DATA_20,
    output  wire    [8:0]   ADC48_DATA_21,
    output  wire    [8:0]   ADC48_DATA_22,
    output  wire    [8:0]   ADC48_DATA_23,
    output  wire    [8:0]   ADC48_DATA_24,
    output  wire    [8:0]   ADC48_DATA_25,
    output  wire    [8:0]   ADC48_DATA_26,
    output  wire    [8:0]   ADC48_DATA_27,
    output  wire    [8:0]   ADC48_DATA_28,
    output  wire    [8:0]   ADC48_DATA_29,
    output  wire    [8:0]   ADC48_DATA_30,
    output  wire    [8:0]   ADC48_DATA_31,
    output  wire    [8:0]   ADC48_DATA_32,
    output  wire    [8:0]   ADC48_DATA_33,
    output  wire    [8:0]   ADC48_DATA_34,
    output  wire    [8:0]   ADC48_DATA_35,
    output  wire    [8:0]   ADC48_DATA_36,
    output  wire    [8:0]   ADC48_DATA_37,
    output  wire    [8:0]   ADC48_DATA_38,
    output  wire    [8:0]   ADC48_DATA_39,
    output  wire    [8:0]   ADC48_DATA_40,
    output  wire    [8:0]   ADC48_DATA_41,
    output  wire    [8:0]   ADC48_DATA_42,
    output  wire    [8:0]   ADC48_DATA_43,
    output  wire    [8:0]   ADC48_DATA_44,
    output  wire    [8:0]   ADC48_DATA_45,
    output  wire    [8:0]   ADC48_DATA_46,
    output  wire    [8:0]   ADC48_DATA_47
);

    reg clk500m;
    reg clk200m;

    // generate clock: T1 = 2ns, T2 = 5ns
    initial begin
        clk500m = 0;
        forever
        begin
            #1 clk500m = ~clk500m;
        end
    end

    initial begin
        clk200m = 0;
        forever
        begin
            #2.5 clk200m = ~clk200m;
        end
    end

    assign CLK500M = clk500m;
    assign CLK200M = clk200m;

endmodule
