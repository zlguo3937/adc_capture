**** Created by MC2: Version 2012.02.00.d on 2024/05/13, 17:41:28 

************************************************************************
* AUCDL NETLIST:
* 
* LIBRARY NAME:  N28HP_SP_LEAFCELLS
* TOP CELL NAME: LEAFCELLS_DR
* VIEW NAME:     SCHEMATIC
* NETLISTED ON:  JAN 18 15:09:47 2013
************************************************************************

*.EQUATION
*.SCALE METER
.PARAM


*.PIN VSS

************************************************************************
* LIBRARY NAME: N28_LOGIC_MAC
* CELL NAME:    NOR_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_NOR_BULK A B G GB P PB Y
*.PININFO A:I B:I G:I GB:I P:I PB:I Y:O
M1 NET021 A P PB pch_mac L=LP1 W=WP1 M=MULTI*FP1
M3 Y B NET021 PB pch_mac L=LP2 W=WP2 M=MULTI*FP2
M5 Y B G GB nch_mac L=LN2 W=WN2 M=MULTI*FN2
M7 Y A G GB nch_mac L=LN1 W=WN1 M=MULTI*FN1
.ENDS

************************************************************************
* LIBRARY NAME: N28_LOGIC_MAC
* CELL NAME:    INV_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_INV_BULK A G GB P PB Y
*.PININFO A:I G:I GB:I P:I PB:I Y:O
M1 Y A P PB pch_mac L=LP W=WP M=MULTI*FP
M3 Y A G GB nch_mac L=LN W=WN M=MULTI*FN
.ENDS

************************************************************************
* LIBRARY NAME: N28_LOGIC_MAC
* CELL NAME:    NAND_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_NAND_BULK A B G GB P PB Y
*.PININFO A:I B:I G:I GB:I P:I PB:I Y:O
M1 Y A P PB pch_mac L=LP1 W=WP1 M=MULTI*FP1
M4 Y B P PB pch_mac L=LP2 W=WP2 M=MULTI*FP2
M6 Y B NET9 GB nch_mac L=LN2 W=WN2 M=MULTI*FN2
M8 NET9 A G GB nch_mac L=LN1 W=WN1 M=MULTI*FN1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    DOUT
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_DOUT AWT AWTD GBL GBLB Q SLP_Q VDDF VDDFHD VDDHD VDDI VSSI WLP_SAEB
*.PININFO AWT:I AWTD:I SLP_Q:I WLP_SAEB:I Q:O GBL:B GBLB:B VDDF:B VDDFHD:B 
*.PININFO VDDHD:B VDDI:B VSSI:B
XI163 AWTB DLRSB VSSI VSSI VDDHD VDDI DSLRP S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.4U 
+ LN1=0.03U FN2=1 WN2=0.4U LN2=0.03U FP2=1 WP2=0.4U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.4U LP1=0.03U
MM15 QB QBB NET085 VDDI pch_mac L=30N W=0.375U M=8
MM7 NET0102 DSLRP VDDHD VDDI pch_mac L=30N W=1U M=2
MM6 NET0101 DSLRP VDDHD VDDI pch_mac L=30N W=1U M=2
MM4 IOBL GBL NET0101 VDDI pch_mac L=30N W=0.5U M=4
MM22 IOBL AWTB NET0136 VDDI pch_mac L=30N W=0.5U M=2
MM20 NET084 QB VDDHD VDDI pch_mac L=30N W=0.5U M=2
MM23 NET0136 AWTD VDDHD VDDI pch_mac L=30N W=0.5U M=2
MM24 IOBLB AWTB NET0128 VDDI pch_mac L=30N W=0.5U M=2
MM5 IOBLB GBLB NET0102 VDDI pch_mac L=30N W=0.5U M=4
MM25 NET0128 AWTDB VDDHD VDDI pch_mac L=30N W=0.5U M=2
MM19 QBB IOBL NET084 VDDI pch_mac L=30N W=0.25U M=4
MP8_MIXV_SLS GBL DLRSB VDDHD VDDI pch_mac L=30N W=0.9U M=5
MP7_MIXV_SLS VDDHD DLRSB GBLB VDDI pch_mac L=30N W=0.9U M=5
MP6 VDDHD GBLB GBL VDDI pch_mac L=30N W=120N M=1
MP0 GBLB GBL VDDHD VDDI pch_mac L=30N W=120N M=1
MM16 NET085 IOBLB VDDHD VDDI pch_mac L=30N W=0.75U M=4
MM12 Q SLP_Q VSSI VSSI nch_mac L=30N W=400N M=1
MM14 QB QBB VSSI VSSI nch_mac L=30N W=250N M=1
MM13 QB IOBLB VSSI VSSI nch_mac L=30N W=0.25U M=4
MM11 IOBLB DSLRN VSSI VSSI nch_mac L=30N W=250N M=1
MM10 IOBLB IOBL VSSI VSSI nch_mac L=30N W=120N M=1
MM9 IOBL IOBLB VSSI VSSI nch_mac L=30N W=120N M=1
MM8 IOBL DSLRN VSSI VSSI nch_mac L=30N W=250N M=1
MM27 IOBLB SLP_Q VSSI VSSI nch_mac L=30N W=200N M=1
MM26 QBB SLP_Q VSSI VSSI nch_mac L=30N W=400N M=1
MM18 QBB QB VSSI VSSI nch_mac L=30N W=250N M=1
MM17 QBB IOBL VSSI VSSI nch_mac L=30N W=0.25U M=4
XI166 AWTD VSSI VSSI VDDHD VDDI AWTDB S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U LN=0.03U MULTI=1 
+ FP=1 WP=0.4U LP=0.03U
XI162 QB VSSI VSSI VDDFHD VDDF Q S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.8U LN=0.03U MULTI=1 FP=4 
+ WP=0.4U LP=0.03U
XI165 AWT VSSI VSSI VDDHD VDDI AWTB S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U LN=0.03U MULTI=1 
+ FP=1 WP=0.4U LP=0.03U
XI160 WLP_SAEB VSSI VSSI VDDHD VDDI DLRSB S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U LN=0.03U 
+ MULTI=1 FP=1 WP=0.4U LP=0.03U
XI164 DLRSB AWT VSSI VSSI VDDHD VDDI DSLRN S1BSVTSWSO8000Y24_NOR_BULK FN1=1 WN1=0.4U LN1=0.03U 
+ FN2=1 WN2=0.4U LN2=0.03U FP2=1 WP2=0.4U LP2=0.03U MULTI=1 FP1=1 WP1=0.4U 
+ LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    DIN_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_DIN_WOBIST AWTD BWEB BWEBM CKD D DM GW GWB SLP_Q VDDHD VDDI VSSI
*.PININFO BWEB:I BWEBM:I CKD:I D:I DM:I SLP_Q:I AWTD:O GW:O GWB:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
XI339 BX4L SLP_Q VSSI VSSI VDDHD VDDI BX4L1B S1BSVTSWSO8000Y24_NOR_BULK FN1=1 WN1=0.27U 
+ LN1=0.03U FN2=1 WN2=0.27U LN2=0.03U FP2=1 WP2=0.52U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.52U LP1=0.03U
MP1 DX4L3B_AND CKD2 VDDI VDDI pch_mac L=30N W=350N M=1
MM27 DX4L DX4 Z9 VDDI pch_mac L=30N W=200N M=1
MM40 BX4L CKD1B Z16 VDDI pch_mac L=30N W=200N M=1
MM39 VDDHD BX4L1B Z16 VDDI pch_mac L=30N W=200N M=1
MM38 VDDHD CKD2 Z13 VDDI pch_mac L=30N W=200N M=1
MM26 VDDHD CKD2 Z9 VDDI pch_mac L=30N W=200N M=1
MM54 DX4L3B_AND BX4L1B VDDI VDDI pch_mac L=30N W=350N M=1
MM53 DX4L2_AND BX4L1B VDDI VDDI pch_mac L=30N W=350N M=1
MM52 DX4L2_AND DX4L1B VDDI VDDI pch_mac L=30N W=350N M=1
MM51 DX4L3B_AND DX4L2 VDDI VDDI pch_mac L=30N W=350N M=1
MP10 DX4L2_AND CKD2 VDDI VDDI pch_mac L=30N W=350N M=1
MM28 VDDHD DX4L1B Z6 VDDI pch_mac L=30N W=200N M=1
MP5 AWTD DX4 Z19 VDDI pch_mac L=30N W=270N M=1
MP4 Z19 BX1B VDDHD VDDI pch_mac L=30N W=270N M=1
MP3 Z18 BX4 VDDHD VDDI pch_mac L=30N W=270N M=1
MP2 AWTD DX1B Z18 VDDI pch_mac L=30N W=270N M=1
MM41 BX4L BX4 Z13 VDDI pch_mac L=30N W=200N M=1
MM29 DX4L CKD1B Z6 VDDI pch_mac L=30N W=200N M=1
MN6 AWTD DX1B Z20 VSSI nch_mac L=30N W=135N M=1
MN13 Z20 DX4 VSSI VSSI nch_mac L=30N W=135N M=1
MM42 BX4L BX4 Z15 VSSI nch_mac L=30N W=120N M=1
MM43 VSSI CKD1B Z15 VSSI nch_mac L=30N W=120N M=1
MM37 VSSI DX4L1B Z7 VSSI nch_mac L=30N W=120N M=1
MN2 Z2 CKD2 Z1 VSSI nch_mac L=30N W=750N M=2
MM34 DX4L DX4 Z11 VSSI nch_mac L=30N W=120N M=1
MM36 VSSI CKD1B Z11 VSSI nch_mac L=30N W=120N M=1
MN33 DX4L3B_AND DX4L2 Z2 VSSI nch_mac L=30N W=375N M=2
MM35 DX4L CKD2 Z7 VSSI nch_mac L=30N W=120N M=1
MN1 DX4L2_AND DX4L1B Z2 VSSI nch_mac L=30N W=375N M=2
MN7 Z1 BX4L1B VSSI VSSI nch_mac L=30N W=750N M=4
MM45 BX4L CKD2 Z14 VSSI nch_mac L=30N W=120N M=1
MM44 VSSI BX4L1B Z14 VSSI nch_mac L=30N W=120N M=1
MN4 Z20 BX1B VSSI VSSI nch_mac L=30N W=135N M=1
MN5 AWTD BX4 Z20 VSSI nch_mac L=30N W=135N M=1
XI331 DX4L1B VSSI VSSI VDDHD VDDI DX4L2 S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.135U LN=0.03U 
+ MULTI=1 FP=1 WP=0.54U LP=0.03U
XI314 CKD VSSI VSSI VDDHD VDDI CKD1B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.14U LN=0.03U MULTI=1 
+ FP=1 WP=0.2U LP=0.03U
XI317 CKD1B VSSI VSSI VDDHD VDDI CKD2 S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.19U LN=0.03U 
+ MULTI=1 FP=2 WP=0.27U LP=0.03U
XI329 DX4L VSSI VSSI VDDHD VDDI DX4L1B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.27U LN=0.03U 
+ MULTI=1 FP=1 WP=0.54U LP=0.03U
XI326 BX1B VSSI VSSI VDDHD VDDI BX4 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.12U LP=0.03U
XI322 DX1B VSSI VSSI VDDHD VDDI DX4 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.12U LP=0.03U
XI333 DX4L3B_AND VSSI VSSI VDDHD VDDI GW S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.15U LN=0.03U 
+ MULTI=1 FP=10 WP=0.45U LP=0.03U
XI325 BWEB VSSI VSSI VDDHD VDDI BX1B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.12U LP=0.03U
XI321 D VSSI VSSI VDDHD VDDI DX1B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.12U LP=0.03U
XI332 DX4L2_AND VSSI VSSI VDDHD VDDI GWB S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.15U LN=0.03U 
+ MULTI=1 FP=10 WP=0.45U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    IO_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_IO_WOBIST AWT BWEB BWEBM CKD D DM GBL GBLB GW GWB Q SLP_Q VDDF VDDFHD 
+ VDDHD VDDI VSSI WLP_SAEB
*.PININFO AWT:I BWEB:I BWEBM:I CKD:I D:I DM:I SLP_Q:I WLP_SAEB:I GW:O GWB:O 
*.PININFO Q:O GBL:B GBLB:B VDDF:B VDDFHD:B VDDHD:B VDDI:B VSSI:B
XDOUT AWT AWTD GBL GBLB Q SLP_Q VDDF VDDFHD VDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_DOUT
XDIN AWTD BWEB BWEBM CKD D DM GW GWB SLP_Q VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DIN_WOBIST
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    IO_M16_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_IO_M16_WOBIST AWT BWEB BWEBM CKD D DM GBL GBLB GW GWB IOPD PDI PDO Q 
+ SLP_Q VDDF VDDFHD VDDHD VDDI VSSI WLP_SAEB
*.PININFO AWT:I BWEB:I BWEBM:I CKD:I D:I DM:I IOPD:I PDI:I SLP_Q:I WLP_SAEB:I 
*.PININFO GW:O GWB:O PDO:O Q:O GBL:B GBLB:B VDDF:B VDDFHD:B VDDHD:B VDDI:B 
*.PININFO VSSI:B
XI1_MIXV_SLS PDI IOPD VSSI VSSI VDDI VDDI NET45 S1BSVTSWSO8000Y24_NOR_BULK FN1=1 WN1=0.5U 
+ LN1=0.035U FN2=1 WN2=0.5U LN2=0.035U FP2=1 WP2=1U LP2=0.035U MULTI=1 FP1=1 
+ WP1=1U LP1=0.035U
MP1 VDDHD PDO VDDI VDDI pch_mac L=35.0N W=1U M=20
XI159_MIXV_SLS NET45 VSSI VSSI VDDI VDDI PDO S1BSVTSWSO8000Y24_INV_BULK FN=8 WN=0.5U LN=0.035U 
+ MULTI=1 FP=8 WP=1U LP=0.035U
XIO AWT BWEB BWEBM CKD D DM GBL GBLB GW GWB Q SLP_Q VDDF VDDFHD VDDHD VDDI 
+ VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_WOBIST
.ENDS

************************************************************************
* LIBRARY NAME: N28_LOGIC_MAC
* CELL NAME:    TRI_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_TRI_BULK A G GB P PB SEL SELB Y
*.PININFO A:I G:I GB:I P:I PB:I SEL:I SELB:I Y:O
M1 NET016 SELB P PB pch_mac L=LP W=WP M=MULTI*FP
MP0 Y A NET016 PB pch_mac L=LP W=WP M=MULTI*FP
M3 NET7 SEL G GB nch_mac L=LN W=WN M=MULTI*FN
MN0 Y A NET7 GB nch_mac L=LN W=WN M=MULTI*FN
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    LCTRL_PM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_LCTRL_PM DSLP_BUF LIOPD SLP_LCTRL VDDI VSSI
*.PININFO DSLP_BUF:I SLP_LCTRL:I LIOPD:O VDDI:B VSSI:B
MM0 NET087 DSLP_BUFB VDDI VDDI pch_mac L=30N W=0.5U M=2
MM1 NET087 NET77 VSSI VSSI nch_mac L=30N W=500N M=1
XI251 CTRLB VSSI VSSI VDDI VDDI CTRL S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.3U LN=0.03U MULTI=1 
+ FP=2 WP=0.6U LP=0.03U
XI232 DSLP_BUFB VSSI VSSI VDDI VDDI LIOPD S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.3U LN=0.03U 
+ MULTI=1 FP=2 WP=0.6U LP=0.03U
XI230 NET087 VSSI VSSI VDDI VDDI NET97 S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.3U LN=0.03U 
+ MULTI=1 FP=2 WP=0.6U LP=0.03U
XI233 DSLP_BUF VSSI VSSI VDDI VDDI DSLP_BUFB S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.3U LN=0.03U 
+ MULTI=1 FP=1 WP=0.6U LP=0.03U
XI234 SLP_LCTRL DSLP_BUF VSSI VSSI VDDI VDDI NET77 S1BSVTSWSO8000Y24_NOR_BULK FN1=1 WN1=0.3U 
+ LN1=0.03U FN2=1 WN2=0.3U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.3U LP1=0.03U
XI250 SLP_LCTRL DSLP_BUFB VSSI VSSI VDDI VDDI CTRLB S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.3U 
+ LN1=0.03U FN2=1 WN2=0.3U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.3U LP1=0.03U
XI237 NET97 VSSI VSSI VDDI VDDI CTRL CTRLB NET087 S1BSVTSWSO8000Y24_TRI_BULK FN=1 WN=0.12U 
+ LN=0.03U MULTI=1 FP=1 WP=0.12U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    XDRV_READ
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_XDRV_READ BS PD_BUF SAEB VDDHD VDDI VSSI WLP_SAE
*.PININFO BS:I PD_BUF:I WLP_SAE:I SAEB:O VDDHD:B VDDI:B VSSI:B
XNAND0_MIXV_SLH BS WLP_SAE VSSI VSSI VDDHD VDDI BS_WLPSAEB S1BSVTSWSO8000Y24_NAND_BULK FN1=3 
+ WN1=1U LN1=0.03U FN2=3 WN2=1U LN2=0.03U FP2=2 WP2=0.75U LP2=0.03U MULTI=1 
+ FP1=2 WP1=0.75U LP1=0.03U
XI426_MIXV_SLH BS_WLPSAEB VSSI VSSI VDDHD VDDI SAEB S1BSVTSWSO8000Y24_INV_BULK FN=4 WN=0.9U 
+ LN=0.03U MULTI=1 FP=7 WP=1U LP=0.03U
MN1_MIXV_SLH SAEB PD_BUF VSSI VSSI nch_mac L=30N W=120N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    XDRV_Y10
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_XDRV_Y10 PD_BUF VDDHD VDDI VSSI WLPY YIN[0] YIN[1] YOUT[0] YOUT[1]
*.PININFO PD_BUF:I WLPY:I YIN[0]:I YIN[1]:I YOUT[0]:O YOUT[1]:O VDDHD:B VDDI:B 
*.PININFO VSSI:B
MM8 MWL2[1] WLPY VDDHD VDDI pch_mac L=30N W=1U M=1
MM6 YOUT[1] MWL2[1] VDDHD VDDI pch_mac L=30N W=1U M=11
MP31 SHARE WLPY VDDHD VDDI pch_mac L=30N W=150N M=2
MM3 MWL2[0] WLPY VDDHD VDDI pch_mac L=30N W=1U M=1
MM1 MWL2[0] YIN[0] VDDHD VDDI pch_mac L=30N W=1U M=1
MM9 MWL2[1] YIN[1] VDDHD VDDI pch_mac L=30N W=1U M=1
MM4 YOUT[0] MWL2[0] VDDHD VDDI pch_mac L=30N W=1U M=11
MN21 SHARE WLPY VSSI VSSI nch_mac L=30N W=1U M=2
MM2 MWL2[0] YIN[0] SHARE VSSI nch_mac L=30N W=1U M=1
MM0 YOUT[1] PD_BUF VSSI VSSI nch_mac L=30N W=120N M=1
MN3 YOUT[0] PD_BUF VSSI VSSI nch_mac L=30N W=120N M=1
MM5 YOUT[0] MWL2[0] VSSI VSSI nch_mac L=30N W=1U M=5
MM7 YOUT[1] MWL2[1] VSSI VSSI nch_mac L=30N W=1U M=5
MM10 MWL2[1] YIN[1] SHARE VSSI nch_mac L=30N W=1U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    XDRV_Y4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_XDRV_Y4 PD_BUF VDDHD VDDI VSSI WLPY YIN[0] YIN[1] YIN[2] YIN[3] 
+ YOUT[0] YOUT[1] YOUT[2] YOUT[3]
*.PININFO PD_BUF:I WLPY:I YIN[0]:I YIN[1]:I YIN[2]:I YIN[3]:I YOUT[0]:O 
*.PININFO YOUT[1]:O YOUT[2]:O YOUT[3]:O VDDHD:B VDDI:B VSSI:B
MM34 YOUT[3] MWL2[3] VSSI VSSI nch_mac L=30N W=0.73U M=8
MM31 MWL2[3] YIN[3] SHARE VSSI nch_mac L=30N W=0.72U M=4
MM29 YOUT[2] PD_BUF VSSI VSSI nch_mac L=30N W=120N M=1
MM28 MWL2[2] YIN[2] SHARE VSSI nch_mac L=30N W=0.72U M=4
MM23 YOUT[1] MWL2[1] VSSI VSSI nch_mac L=30N W=0.73U M=8
MM19 YOUT[1] PD_BUF VSSI VSSI nch_mac L=30N W=120N M=1
MM26 YOUT[2] MWL2[2] VSSI VSSI nch_mac L=30N W=0.73U M=8
MN3 YOUT[0] PD_BUF VSSI VSSI nch_mac L=30N W=120N M=1
MM36 YOUT[3] PD_BUF VSSI VSSI nch_mac L=30N W=120N M=1
MM2 MWL2[0] YIN[0] SHARE VSSI nch_mac L=30N W=0.72U M=4
MM5 YOUT[0] MWL2[0] VSSI VSSI nch_mac L=30N W=0.73U M=8
MN21 SHARE WLPY VSSI VSSI nch_mac L=30N W=0.8U M=8
MM21 MWL2[1] YIN[1] SHARE VSSI nch_mac L=30N W=0.72U M=4
MM1 MWL2[0] YIN[0] VDDHD VDDI pch_mac L=30N W=0.68U M=3
MM24 YOUT[1] MWL2[1] VDDHD VDDI pch_mac L=30N W=0.8U M=14
MM3 MWL2[0] WLPY VDDHD VDDI pch_mac L=30N W=0.68U M=3
MM25 YOUT[2] MWL2[2] VDDHD VDDI pch_mac L=30N W=0.8U M=14
MP31 SHARE WLPY VDDHD VDDI pch_mac L=30N W=150N M=2
MM4 YOUT[0] MWL2[0] VDDHD VDDI pch_mac L=30N W=0.8U M=14
MM32 MWL2[3] YIN[3] VDDHD VDDI pch_mac L=30N W=0.68U M=3
MM30 MWL2[2] WLPY VDDHD VDDI pch_mac L=30N W=0.68U M=3
MM20 MWL2[1] WLPY VDDHD VDDI pch_mac L=30N W=0.68U M=3
MM33 MWL2[3] WLPY VDDHD VDDI pch_mac L=30N W=0.68U M=3
MM35 YOUT[3] MWL2[3] VDDHD VDDI pch_mac L=30N W=0.8U M=14
MM27 MWL2[2] YIN[2] VDDHD VDDI pch_mac L=30N W=0.68U M=3
MM22 MWL2[1] YIN[1] VDDHD VDDI pch_mac L=30N W=0.68U M=3
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    LCTRL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_LCTRL BLEQB_DN BLEQB_UP DEC_X3_DN DEC_X3_UP DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RE_LIO SAEB VDDHD VDDI VSSI WE WE_LIO 
+ WLP_SAE YL[0] YL[1] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQB_DN:I BLEQB_UP:I DEC_X3_DN:I DEC_X3_UP:I DEC_Y[0]:I DEC_Y[1]:I 
*.PININFO DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I DEC_Y[6]:I DEC_Y[7]:I 
*.PININFO PD_BUF:I RE:I WE:I WLP_SAE:I YL[0]:I YL[1]:I DEC_Y_DN[0]:O 
*.PININFO DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O DEC_Y_DN[4]:O 
*.PININFO DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O DEC_Y_UP[0]:O 
*.PININFO DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O DEC_Y_UP[4]:O 
*.PININFO DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE_LIO:O SAEB:O WE_LIO:O 
*.PININFO YL_LIO[0]:O YL_LIO[1]:O VDDHD:B VDDI:B VSSI:B
XNOR0_MIXV_SSH DEC_X3_UP DEC_X3_DN VSSI VSSI VDDHD VDDI BS0 S1BSVTSWSO8000Y24_NOR_BULK FN1=1 
+ WN1=0.4U LN1=0.03U FN2=1 WN2=0.4U LN2=0.03U FP2=1 WP2=0.5U LP2=0.03U MULTI=1 
+ FP1=1 WP1=0.5U LP1=0.03U
XNAND0_MIXV_SSH BS0 BS5 VSSI VSSI VDDHD VDDI BSD S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.3U 
+ LN1=0.03U FN2=1 WN2=0.3U LN2=0.03U FP2=1 WP2=0.75U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.75U LP1=0.03U
XXDRV_READ BSD PD_BUF SAEB VDDHD VDDI VSSI WLP_SAE S1BSVTSWSO8000Y24_XDRV_READ
XXDRV_RW PD_BUF VDDHD VDDI VSSI BSD RE WE RE_LIO WE_LIO S1BSVTSWSO8000Y24_XDRV_Y10
XXDRV_YL PD_BUF VDDHD VDDI VSSI BSD YL[0] YL[1] YL_LIO[0] YL_LIO[1] S1BSVTSWSO8000Y24_XDRV_Y10
XINV4_MIXV_SSH BS4 VSSI VSSI VDDHD VDDI BS4B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV5_MIXV_SSH BS4B VSSI VSSI VDDHD VDDI BS5 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV0_MIXV_SSH BS0 VSSI VSSI VDDHD VDDI BS1B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV3_MIXV_SSH BS3B VSSI VSSI VDDHD VDDI BS4 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV2_MIXV_SSH BS2 VSSI VSSI VDDHD VDDI BS3B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV1_MIXV_SSH BS1B VSSI VSSI VDDHD VDDI BS2 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XXDRV_Y4_D[0] PD_BUF VDDHD VDDI VSSI BLEQB_DN DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] S1BSVTSWSO8000Y24_XDRV_Y4
XXDRV_Y4_D[1] PD_BUF VDDHD VDDI VSSI BLEQB_DN DEC_Y[4] DEC_Y[5] DEC_Y[6] 
+ DEC_Y[7] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] S1BSVTSWSO8000Y24_XDRV_Y4
XXDRV_Y4_U[0] PD_BUF VDDHD VDDI VSSI BLEQB_UP DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] S1BSVTSWSO8000Y24_XDRV_Y4
XXDRV_Y4_U[1] PD_BUF VDDHD VDDI VSSI BLEQB_UP DEC_Y[4] DEC_Y[5] DEC_Y[6] 
+ DEC_Y[7] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] S1BSVTSWSO8000Y24_XDRV_Y4
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    XDRV_LA512_SHA
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_XDRV_LA512_SHA DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD SLP_LCTRL TK VDDHD VDDI VSSI WE 
+ WLOUT[0] WLOUT[1] WLPY WLPYB WLP_SAE WLP_SAE_TK YL[0] YL[1]
*.PININFO DSLP_BUF:I SLP_LCTRL:I WLPY:I WLPYB:I WLP_SAE:I WLOUT[0]:O 
*.PININFO WLOUT[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B RE:B SH_NPD:B TK:B VDDHD:B VDDI:B VSSI:B WE:B 
*.PININFO WLP_SAE_TK:B YL[0]:B YL[1]:B
MP20_MIXV_SLH WLOUT[0] MWL2 VDDHD VDDI pch_mac L=35.0N W=0.875U M=6
MP4 VDDHD SLP_LCTRL VDDI VDDI pch_mac L=35.0N W=0.75U M=4
MP7 MWL0 DEC_X1[0] VDDI VDDI pch_mac L=35.0N W=100N M=1
MP14 MWL0A DEC_X0[1] VDDI VDDI pch_mac L=35.0N W=100N M=1
MM1_MIXV_SLH WLOUT[1] MWL2A VDDHD VDDI pch_mac L=35.0N W=0.875U M=6
MM3 VDDI WLPY MWL2A VDDI pch_mac L=35.0N W=0.64U M=2
MM8 MWL2 MWL1 VDDI VDDI pch_mac L=35.0N W=0.5U M=2
MM5 MWL2A MWL1A VDDI VDDI pch_mac L=35.0N W=0.5U M=2
MP19 VDDI WLPY MWL2 VDDI pch_mac L=35.0N W=0.64U M=2
MP13 MWL0A DEC_X1[0] VDDI VDDI pch_mac L=35.0N W=100N M=1
MP6 MWL0 DEC_X0[0] VDDI VDDI pch_mac L=35.0N W=100N M=1
MN7 MWL0A DEC_X0[1] SH_NPD VSSI nch_mac L=35.0N W=100N M=1
MN0 MWL2 MWL1 WLPYB VSSI nch_mac L=35.0N W=0.9U M=2
MP9 MWL0 DEC_X0[0] SH_NPD VSSI nch_mac L=35.0N W=100N M=1
MM2_MIXV_SLH WLOUT[1] MWL2A VSSI VSSI nch_mac L=35.0N W=0.65U M=4
MM4 MWL2A MWL1A WLPYB VSSI nch_mac L=35.0N W=0.9U M=2
MN6_MIXV_SLH WLOUT[0] MWL2 VSSI VSSI nch_mac L=35.0N W=0.65U M=4
XI426 MWL0A VSSI VSSI VDDHD VDDI MWL1A S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.39U LN=0.03U 
+ MULTI=1 FP=1 WP=0.565U LP=0.03U
XI425 MWL0 VSSI VSSI VDDHD VDDI MWL1 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.39U LN=0.03U MULTI=1 
+ FP=1 WP=0.565U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    TKBL_EDGE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_TKBL_EDGE BLB_EDGE BL_EDGE G_FLOAT VDDAI VDDI VSSI WL WL_TK TIEH
*.PININFO WL:I WL_TK:I BLB_EDGE:B BL_EDGE:B G_FLOAT:B VDDAI:B VDDI:B VSSI:B 
*.PININFO TIEH:B
MPCHPU1 BLB TIEH VDDAI VDDI pchpu_sr L=35N W=40N M=1
MPCHPU0 VDDAI BLB TIEH VDDI pchpu_sr L=35N W=40N M=1
MNCHPD1 BLB TIEH VSSI VSSI nchpd_sr L=35N W=95N M=1
MNCHPD0 G_FLOAT BLB TIEH VSSI nchpd_sr L=35N W=95N M=1
MNCHPG1 BLB WL BL_EDGE VSSI nchpg_sr L=35N W=65N M=1
MNCHPG0 BLB_EDGE WL TIEH VSSI nchpg_sr L=35N W=65N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28_LOGIC_MAC
* CELL NAME:    AINV
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_AINV A G V Y
*.PININFO A:I G:I V:I Y:O
M1 Y A V V pch_mac L=LP W=WP M=MULTI*FP
M3 Y A G G nch_mac L=LN W=WN M=MULTI*FN
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    DECB1_BS_SEG
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_DECB1_BS_SEG CKP CLK DEC EN ENC PREDEC VDDHD VDDI VSSI
*.PININFO CKP:I CLK:I EN:I ENC:I PREDEC:I DEC:O VDDHD:B VDDI:B VSSI:B
MM3 NT1 PREDEC VDDHD VDDI pch_mac L=30N W=400N M=1
MP5 NT1 EN VDDHD VDDI pch_mac L=30N W=400N M=2
MM2 NT1 CKP NET59 VDDI pch_mac L=30N W=400N M=1
MP0 DEC NT1 VDDHD VDDI pch_mac L=30N W=0.6U M=14
MM1 NET59 CLK VDDHD VDDI pch_mac L=30N W=400N M=1
MTN1 NT1 CKP NT3 VSSI nch_mac L=30N W=400N M=1
MTN2 NT3 PREDEC ENC VSSI nch_mac L=30N W=0.6U M=4
MM0 NT1 CLK NT3 VSSI nch_mac L=30N W=0.6U M=2
MN0 DEC NT1 VSSI VSSI nch_mac L=30N W=0.6U M=7
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    DECB1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_DECB1 CKP CLK DEC EN ENC PREDEC VDDHD VDDI VSSI
*.PININFO CKP:I CLK:I EN:I ENC:I PREDEC:I DEC:O VDDHD:B VDDI:B VSSI:B
MTN1 NT1 CKP NT3 VSSI nch_mac L=30N W=400N M=1
MTN2 NT3 PREDEC ENC VSSI nch_mac L=30N W=0.6U M=4
MM0 NT1 CLK NT3 VSSI nch_mac L=30N W=0.6U M=2
MN0 DEC NT1 VSSI VSSI nch_mac L=30N W=0.6U M=7
MM1 NET65 CLK VDDHD VDDI pch_mac L=30N W=400N M=1
MM3 NT1 PREDEC VDDHD VDDI pch_mac L=30N W=400N M=1
MP0 DEC NT1 VDDHD VDDI pch_mac L=30N W=0.6U M=14
MP5 NT1 EN VDDHD VDDI pch_mac L=30N W=400N M=2
MM2 NT1 CKP NET65 VDDI pch_mac L=30N W=400N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    DECB4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_DECB4 IN0A IN0B IN1A IN1B IN2 PREDEC0 PREDEC1 PREDEC2 PREDEC3 VDDHD 
+ VDDI VSSI
*.PININFO IN0A:I IN0B:I IN1A:I IN1B:I IN2:I PREDEC0:O PREDEC1:O PREDEC2:O 
*.PININFO PREDEC3:O VDDHD:B VDDI:B VSSI:B
MM19 N5 IN1B NET19 VSSI nch_mac L=30N W=420N M=1
MM20 NET0154 IN0B N5 VSSI nch_mac L=30N W=195N M=1
MM21 NET0150 IN0A N5 VSSI nch_mac L=30N W=195N M=1
MM26 NET19 IN2 VSSI VSSI nch_mac L=30N W=420N M=2
MM8 N2 IN1A NET19 VSSI nch_mac L=30N W=420N M=1
MM7 NET0138 IN0B N2 VSSI nch_mac L=30N W=195N M=1
MM0 NET0134 IN0A N2 VSSI nch_mac L=30N W=195N M=1
MM15 NET0154 IN1B VDDHD VDDI pch_mac L=30N W=200N M=1
MM16 NET0154 IN0B VDDHD VDDI pch_mac L=30N W=200N M=1
MM17 NET0150 IN1B VDDHD VDDI pch_mac L=30N W=200N M=1
MM18 NET0150 IN0A VDDHD VDDI pch_mac L=30N W=200N M=1
MM22 NET0150 IN2 VDDHD VDDI pch_mac L=30N W=200N M=1
MM23 NET0154 IN2 VDDHD VDDI pch_mac L=30N W=200N M=1
MM24 NET0138 IN2 VDDHD VDDI pch_mac L=30N W=200N M=1
MM25 NET0134 IN2 VDDHD VDDI pch_mac L=30N W=200N M=1
MM5 NET0138 IN1A VDDHD VDDI pch_mac L=30N W=200N M=1
MM4 NET0138 IN0B VDDHD VDDI pch_mac L=30N W=200N M=1
MM2 NET0134 IN1A VDDHD VDDI pch_mac L=30N W=200N M=1
MM1 NET0134 IN0A VDDHD VDDI pch_mac L=30N W=200N M=1
XINV3 NET0154 VSSI VSSI VDDHD VDDI PREDEC3 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.195U LN=0.03U 
+ MULTI=1 FP=2 WP=0.2U LP=0.03U
XINV2 NET0150 VSSI VSSI VDDHD VDDI PREDEC2 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.195U LN=0.03U 
+ MULTI=1 FP=2 WP=0.2U LP=0.03U
XINV1 NET0138 VSSI VSSI VDDHD VDDI PREDEC1 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.195U LN=0.03U 
+ MULTI=1 FP=2 WP=0.2U LP=0.03U
XINV0 NET0134 VSSI VSSI VDDHD VDDI PREDEC0 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.195U LN=0.03U 
+ MULTI=1 FP=2 WP=0.2U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    ABUF_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_ABUF_WOBIST A AC AM AXL AX1B BIST1B BIST2 CK1B CK2 VDDHD VDDI VSSI
*.PININFO A:I AM:I BIST1B:I BIST2:I CK1B:I CK2:I AC:O AXL:O AX1B:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
MM23 NET0108 CK1B VSSI VSSI nch_mac L=30N W=750N M=1
MM21 NET078 AC VSSI VSSI nch_mac L=30N W=120N M=1
MM20 AXL CK2 NET078 VSSI nch_mac L=30N W=120N M=1
MM19 AXL A NET0108 VSSI nch_mac L=30N W=750N M=1
MM29 AXL A NET0145 VDDI pch_mac L=30N W=750N M=1
MM28 NET0145 CK2 VDDHD VDDI pch_mac L=30N W=0.75U M=2
MM27 NET0149 AC VDDHD VDDI pch_mac L=30N W=120N M=1
MM26 AXL CK1B NET0149 VDDI pch_mac L=30N W=120N M=1
XI25 AXL VSSI VSSI VDDHD VDDI AC S1BSVTSWSO8000Y24_INV_BULK FN=3 WN=0.2U LN=0.03U MULTI=1 FP=3 
+ WP=0.3U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    ABUF_DECB4_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_ABUF_DECB4_WOBIST AX[0] AX[1] AX[2] BIST1B BIST2 CK1B CK2 IN[0] IN[1] 
+ IN[2] IN_M[0] IN_M[1] IN_M[2] OUT[0] OUT[1] OUT[2] OUT[3] OUT[4] OUT[5] 
+ OUT[6] OUT[7] VDDHD VDDI VSSI
*.PININFO BIST1B:I BIST2:I CK1B:I CK2:I IN[0]:I IN[1]:I IN[2]:I IN_M[0]:I 
*.PININFO IN_M[1]:I IN_M[2]:I AX[0]:O AX[1]:O AX[2]:O OUT[0]:O OUT[1]:O 
*.PININFO OUT[2]:O OUT[3]:O OUT[4]:O OUT[5]:O OUT[6]:O OUT[7]:O VDDHD:B VDDI:B 
*.PININFO VSSI:B
XABUF[0] IN[0] AXC[0] IN_M[0] AXT[0] AX[0] BIST1B BIST2 CK1B CK2 VDDHD VDDI 
+ VSSI S1BSVTSWSO8000Y24_ABUF_WOBIST
XABUF[1] IN[1] AXC[1] IN_M[1] AXT[1] AX[1] BIST1B BIST2 CK1B CK2 VDDHD VDDI 
+ VSSI S1BSVTSWSO8000Y24_ABUF_WOBIST
XABUF[2] IN[2] AXC[2] IN_M[2] AXT[2] AX[2] BIST1B BIST2 CK1B CK2 VDDHD VDDI 
+ VSSI S1BSVTSWSO8000Y24_ABUF_WOBIST
XDECB4[0] AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] OUT[0] OUT[1] OUT[2] OUT[3] VDDHD 
+ VDDI VSSI S1BSVTSWSO8000Y24_DECB4
XDECB4[1] AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] OUT[4] OUT[5] OUT[6] OUT[7] VDDHD 
+ VDDI VSSI S1BSVTSWSO8000Y24_DECB4
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    DECB2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_DECB2 IN0A IN0B IN1 PREDEC0 PREDEC1 VDDHD VDDI VSSI
*.PININFO IN0A:I IN0B:I IN1:I PREDEC0:O PREDEC1:O VDDHD:B VDDI:B VSSI:B
MM0 N1 IN0A N2 VSSI nch_mac L=30N W=195N M=1
MM7 N3 IN0B N2 VSSI nch_mac L=30N W=195N M=1
MM8 N2 IN1 VSSI VSSI nch_mac L=30N W=420N M=1
MM2 N1 IN1 VDDHD VDDI pch_mac L=30N W=200N M=1
MM1 N1 IN0A VDDHD VDDI pch_mac L=30N W=200N M=1
MM5 N3 IN1 VDDHD VDDI pch_mac L=30N W=200N M=1
MM4 N3 IN0B VDDHD VDDI pch_mac L=30N W=200N M=1
XINV0 N3 VSSI VSSI VDDHD VDDI PREDEC1 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.195U LN=0.03U 
+ MULTI=1 FP=2 WP=0.2U LP=0.03U
XINV1 N1 VSSI VSSI VDDHD VDDI PREDEC0 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.195U LN=0.03U 
+ MULTI=1 FP=2 WP=0.2U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    ABUF_DECB2_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_ABUF_DECB2_WOBIST AX[0] AX[1] BIST1B BIST2 CK1B CK2 IN[0] IN[1] 
+ IN_M[0] IN_M[1] OUT[0] OUT[1] OUT[2] OUT[3] VDDHD VDDI VSSI
*.PININFO BIST1B:I BIST2:I CK1B:I CK2:I IN[0]:I IN[1]:I IN_M[0]:I IN_M[1]:I 
*.PININFO AX[0]:O AX[1]:O OUT[0]:O OUT[1]:O OUT[2]:O OUT[3]:O VDDHD:B VDDI:B 
*.PININFO VSSI:B
XABUF[0] IN[0] AXC[0] IN_M[0] AXT[0] AX[0] BIST1B BIST2 CK1B CK2 VDDHD VDDI 
+ VSSI S1BSVTSWSO8000Y24_ABUF_WOBIST
XABUF[1] IN[1] AXC[1] IN_M[1] AXT[1] AX[1] BIST1B BIST2 CK1B CK2 VDDHD VDDI 
+ VSSI S1BSVTSWSO8000Y24_ABUF_WOBIST
XDECB2[0] AXC[0] AXT[0] AXC[1] OUT[0] OUT[1] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB2
XDECB2[1] AXC[0] AXT[0] AXT[1] OUT[2] OUT[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB2
.ENDS

************************************************************************
* LIBRARY NAME: N28_LOGIC_MAC
* CELL NAME:    NAND3_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_NAND3_BULK A B C G GB P PB Y
*.PININFO A:I B:I C:I G:I GB:I P:I PB:I Y:O
M1 Y A P PB pch_mac L=LP1 W=WP1 M=MULTI*FP1
M3 Y B P PB pch_mac L=LP2 W=WP2 M=MULTI*FP2
M7 Y C P PB pch_mac L=LP3 W=WP3 M=MULTI*FP3
M9 Y C NET17 GB nch_mac L=LN3 W=WN3 M=MULTI*FN3
M11 NET17 B NET14 GB nch_mac L=LN2 W=WN2 M=MULTI*FN2
M13 NET14 A G GB nch_mac L=LN1 W=WN1 M=MULTI*FN1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    RESETD_TSEL_WT
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_RESETD_TSEL_WT CKPB TK VDDHD VDDI VSSI OUT WV[0] WV[1]
*.PININFO CKPB:I WV[0]:I WV[1]:I OUT:O TK:B VDDHD:B VDDI:B VSSI:B
XI87_MIXV_SSH TD_01_11 TD_10 VSSI VSSI VDDHD VDDI NET78 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 
+ WN1=0.375U LN1=0.03U FN2=1 WN2=0.375U LN2=0.03U FP2=1 WP2=0.27U LP2=0.03U 
+ MULTI=1 FP1=1 WP1=0.27U LP1=0.03U
XND0_MIXV_SSH CKPB TD_10 VSSI VSSI VDDHD VDDI Z0 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.375U 
+ LN1=0.03U FN2=1 WN2=0.375U LN2=0.03U FP2=1 WP2=0.27U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.27U LP1=0.03U
XND5_MIXV_SSH Z5 WV[1] VSSI VSSI VDDHD VDDI TD_10 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.375U 
+ LN1=0.03U FN2=1 WN2=0.375U LN2=0.03U FP2=1 WP2=0.2U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.2U LP1=0.03U
XI84_MIXV_SSH Z0 WV[0] VSSI VSSI VDDHD VDDI TD_01_11 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 
+ WN1=0.375U LN1=0.03U FN2=1 WN2=0.375U LN2=0.03U FP2=1 WP2=0.27U LP2=0.03U 
+ MULTI=1 FP1=1 WP1=0.27U LP1=0.03U
XI83_MIXV_SSH Z4 VSSI VSSI VDDHD VDDI Z5 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.18U LP=0.03U
XI65_MIXV_SSH Z3 VSSI VSSI VDDHD VDDI Z4 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.18U LP=0.03U
XI64_MIXV_SSH CKPB VSSI VSSI VDDHD VDDI Z3 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.18U LP=0.03U
XI89_MIXV_SSH NET78 VSSI VSSI VDDHD VDDI OUT S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.18U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    PMCTRL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_PMCTRL CKP DSLP DSLP_BUF SD SD_BUF SLP SLP_BUF VDDI VSSI
*.PININFO CKP:I DSLP:I SD:I SLP:I DSLP_BUF:O SD_BUF:O SLP_BUF:O VDDI:B VSSI:B
XI63 NET072 VSSI VDDI SLP_BUF S1BSVTSWSO8000Y24_AINV FN=4 WN=300N LN=0.03U MULTI=1 FP=4 
+ WP=600N LP=0.03U
XI62 NET084 VSSI VDDI DSLP_BUF S1BSVTSWSO8000Y24_AINV FN=4 WN=300N LN=0.03U MULTI=1 FP=4 
+ WP=600N LP=0.03U
XI61 NET088 VSSI VDDI SD_BUF4 S1BSVTSWSO8000Y24_AINV FN=4 WN=300N LN=0.03U MULTI=1 FP=4 
+ WP=600N LP=0.03U
XI68 NET0111 VSSI VDDI SLP_BUF1 S1BSVTSWSO8000Y24_AINV FN=1 WN=300N LN=0.03U MULTI=1 FP=1 
+ WP=600N LP=0.03U
XI66 NET030 VSSI VDDI DSLP_BUF1 S1BSVTSWSO8000Y24_AINV FN=1 WN=300N LN=0.03U MULTI=1 FP=1 
+ WP=600N LP=0.03U
XI53 SD_BUF VSSI VDDI NET088 S1BSVTSWSO8000Y24_AINV FN=1 WN=300N LN=0.03U MULTI=1 FP=1 WP=600N 
+ LP=0.03U
XI57 DSLP_BUF1 VSSI VDDI NET084 S1BSVTSWSO8000Y24_AINV FN=1 WN=300N LN=0.03U MULTI=1 FP=1 
+ WP=600N LP=0.03U
XI48 SD VSSI VDDI NET0129 S1BSVTSWSO8000Y24_AINV FN=1 WN=300N LN=0.03U MULTI=1 FP=1 WP=600N 
+ LP=0.03U
XI60 SLP_BUF1 VSSI VDDI NET072 S1BSVTSWSO8000Y24_AINV FN=1 WN=300N LN=0.03U MULTI=1 FP=1 
+ WP=600N LP=0.03U
XI49 NET0129 VSSI VDDI SD_BUF S1BSVTSWSO8000Y24_AINV FN=1 WN=300N LN=0.03U MULTI=1 FP=1 
+ WP=600N LP=0.03U
XI44 DSLP_BUF1 SLP VSSI VSSI VDDI VDDI NET0111 S1BSVTSWSO8000Y24_NOR_BULK FN1=1 WN1=0.3U 
+ LN1=0.03U FN2=1 WN2=0.3U LN2=0.03U FP2=1 WP2=0.6U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.6U LP1=0.03U
XI37 SD_BUF DSLP VSSI VSSI VDDI VDDI NET030 S1BSVTSWSO8000Y24_NOR_BULK FN1=1 WN1=0.3U 
+ LN1=0.03U FN2=1 WN2=0.3U LN2=0.03U FP2=1 WP2=0.6U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.6U LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    DECB1_DCLK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_DECB1_DCLK CKP CLK DEC EN ENC PREDEC VDDHD VDDI VSSI
*.PININFO CKP:I CLK:I EN:I ENC:I PREDEC:I DEC:O VDDHD:B VDDI:B VSSI:B
MM0 NT1 CLK NT3 VSSI nch_mac L=30N W=0.6U M=2
MN0 DEC NT1 VSSI VSSI nch_mac L=30N W=0.6U M=6
MTN1 NT1 CKP NT3 VSSI nch_mac L=30N W=400N M=1
MTN2 NT3 PREDEC ENC VSSI nch_mac L=30N W=0.6U M=3
MP5 NT1 EN VDDHD VDDI pch_mac L=30N W=400N M=1
MM2 NT1 CKP NET59 VDDI pch_mac L=30N W=400N M=1
MM1 NET59 CLK VDDHD VDDI pch_mac L=30N W=400N M=1
MM3 NT1 PREDEC VDDHD VDDI pch_mac L=30N W=400N M=1
MP0 DEC NT1 VDDHD VDDI pch_mac L=30N W=0.6U M=12
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    CKBUF_M8_DR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_CKBUF_M8_DR CK1B CK2 CKP CLK VDDHD VDDI VSSI
*.PININFO CKP:I CLK:I CK1B:O CK2:O VDDHD:B VDDI:B VSSI:B
XINV0 CK1B VSSI VSSI VDDHD VDDI CK2 S1BSVTSWSO8000Y24_INV_BULK FN=4 WN=0.54U LN=0.03U MULTI=1 
+ FP=4 WP=1U LP=0.03U
XNOR0 CLK CKP VSSI VSSI VDDHD VDDI CK1B S1BSVTSWSO8000Y24_NOR_BULK FN1=2 WN1=0.8U LN1=0.03U 
+ FN2=1 WN2=0.375U LN2=0.03U FP2=3 WP2=1U LP2=0.03U MULTI=1 FP1=3 WP1=1U 
+ LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    ENBUFB_M8_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_ENBUFB_M8_WOBIST BIST1B BIST2 CEBX CEBM CK1B CK2 EN ENC EN_D EN_DCLK 
+ RSC VDDHD VDDI VSSI
*.PININFO BIST1B:I BIST2:I CEBX:I CEBM:I CK1B:I CK2:I RSC:I EN:O ENC:O EN_D:O 
*.PININFO EN_DCLK:O VDDHD:B VDDI:B VSSI:B
XI158 NET109 NET109 VSSI VSSI VDDHD VDDI NET100 S1BSVTSWSO8000Y24_NOR_BULK FN1=1 WN1=0.12U 
+ LN1=0.03U FN2=1 WN2=0.12U LN2=0.03U FP2=1 WP2=0.12U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.12U LP1=0.03U
MN100 ENC EN VSSI VSSI nch_mac L=30N W=1.21U M=1
MM5 NET0188 RSC VSSI VSSI nch_mac L=30N W=270N M=1
MM4 NET0168 EN NET0188 VSSI nch_mac L=30N W=135N M=1
MM3 CEBXL CK2 NET0168 VSSI nch_mac L=30N W=135N M=1
MM20 NET0151 RSC VSSI VSSI nch_mac L=30N W=1.125U M=1
MM17 CEBXL CEBX NET0253 VSSI nch_mac L=30N W=630N M=1
MM18 NET0253 CK1B NET0151 VSSI nch_mac L=30N W=630N M=1
MN300 ENC EN VSSI VSSI nch_mac L=30N W=1.31U M=13
MM19 NET0286 CK2 VDDI VDDI pch_mac L=30N W=1.125U M=1
MM2 NET0203 EN VDDI VDDI pch_mac L=30N W=195N M=1
MM7 CEBXL RSC VDDI VDDI pch_mac L=30N W=750N M=1
MM16 CEBXL CEBX NET0286 VDDI pch_mac L=30N W=1.125U M=1
MM1 CEBXL CK1B NET0203 VDDI pch_mac L=30N W=195N M=1
XINV7 NET0183 VSSI VSSI VDDHD VDDI NET115 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XI147 NET0179 VSSI VSSI VDDHD VDDI NET0183 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XI148 EN VSSI VSSI VDDHD VDDI NET0179 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV8 NET115 VSSI VSSI VDDHD VDDI NET109 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XI152 NET94 VSSI VSSI VDDHD VDDI EN_D S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=1.125U LN=0.03U 
+ MULTI=1 FP=4 WP=1.1U LP=0.03U
XINV5 EN VSSI VSSI VDDI VDDI NET94 S1BSVTSWSO8000Y24_INV_BULK FN=3 WN=0.35U LN=0.03U MULTI=1 
+ FP=1 WP=0.54U LP=0.03U
XI161 EN VSSI VSSI VDDHD VDDI NET0170 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=150N LN=0.03U MULTI=1 
+ FP=1 WP=300N LP=0.03U
XI157 NET0170 VSSI VSSI VDDHD VDDI EN_DCLK S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=300N LN=0.03U 
+ MULTI=1 FP=2 WP=300N LP=0.03U
XI141 CEBXL VSSI VSSI VDDI VDDI EN S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=1.14U LN=0.03U MULTI=1 
+ FP=4 WP=1.125U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    CDEC_M8_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_CDEC_M8_WOBIST AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] 
+ AX[9] AX[10] BIST1B BIST2 CEB CEBM CK2 CKD CKP CKPD CKPDCLK CLK CLK_DR 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN 
+ RE REDEN REDENB RSC VDDHD VDDI VSSI WE WEB WEB3B WEBM X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] 
+ YM[2] YM[3]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CKPDCLK:I CLK:I CLK_DR:I 
*.PININFO REDEN:I REDENB:I RSC:I WEB:I WEBM:I X[0]:I X[1]:I X[2]:I X[3]:I 
*.PININFO X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I 
*.PININFO XM[10]:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I 
*.PININFO AX[0]:O AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O AX[6]:O AX[7]:O 
*.PININFO AX[8]:O AX[9]:O AX[10]:O CK2:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O 
*.PININFO DEC_X3[2]:O DEC_X3[3]:O DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O 
*.PININFO DEC_X3[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O 
*.PININFO DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O EN:O RE:O WE:O WEB3B:O YL[0]:O 
*.PININFO YL[1]:O VDDHD:B VDDI:B VSSI:B
XIDEC_Y[0] CKPD CLK_DR DEC_Y[0] EN_D ENC XY[0] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_Y[1] CKPD CLK_DR DEC_Y[1] EN_D ENC XY[1] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_Y[2] CKPD CLK_DR DEC_Y[2] EN_D ENC XY[2] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_Y[3] CKPD CLK_DR DEC_Y[3] EN_D ENC XY[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_Y[4] CKPD CLK_DR DEC_Y[4] EN_D ENC XY[4] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_Y[5] CKPD CLK_DR DEC_Y[5] EN_D ENC XY[5] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_Y[6] CKPD CLK_DR DEC_Y[6] EN_D ENC XY[6] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_Y[7] CKPD CLK_DR DEC_Y[7] EN_D ENC XY[7] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_WE CKPD CLK_DR WE EN_D ENC WEB3B VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X1[0] CKPD CLK_DR DEC_X1[0] EN_D ENC XB[0] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X1[1] CKPD CLK_DR DEC_X1[1] EN_D ENC XB[1] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X1[2] CKPD CLK_DR DEC_X1[2] EN_D ENC XB[2] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X1[3] CKPD CLK_DR DEC_X1[3] EN_D ENC XB[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X1[4] CKPD CLK_DR DEC_X1[4] EN_D ENC XB[4] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X1[5] CKPD CLK_DR DEC_X1[5] EN_D ENC XB[5] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X1[6] CKPD CLK_DR DEC_X1[6] EN_D ENC XB[6] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X1[7] CKPD CLK_DR DEC_X1[7] EN_D ENC XB[7] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X2[0] CKPD CLK_DR DEC_X2[0] EN_D ENC XC[0] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X2[1] CKPD CLK_DR DEC_X2[1] EN_D ENC XC[1] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X2[2] CKPD CLK_DR DEC_X2[2] EN_D ENC XC[2] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X2[3] CKPD CLK_DR DEC_X2[3] EN_D ENC XC[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_YL[0] CKPD CLK_DR YL[0] EN_D ENC AYC[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_YL[1] CKPD CLK_DR YL[1] EN_D ENC AYC1B[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_RE CKPD CLK_DR RE EN_D ENC WEB4 VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X0[0] CKPD CLK_DR DEC_X0[0] EN_D ENC XA[0] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X0[1] CKPD CLK_DR DEC_X0[1] EN_D ENC XA[1] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X0[2] CKPD CLK_DR DEC_X0[2] EN_D ENC XA[2] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X0[3] CKPD CLK_DR DEC_X0[3] EN_D ENC XA[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X0[4] CKPD CLK_DR DEC_X0[4] EN_D ENC XA[4] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X0[5] CKPD CLK_DR DEC_X0[5] EN_D ENC XA[5] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X0[6] CKPD CLK_DR DEC_X0[6] EN_D ENC XA[6] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XIDEC_X0[7] CKPD CLK_DR DEC_X0[7] EN_D ENC XA[7] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1
XWEBBUF WEB WEB3B WEBM WEB2 WEBX BIST1B BIST2 CK1B CK2 VDDHD VDDI VSSI 
+ S1BSVTSWSO8000Y24_ABUF_WOBIST
XABUF_Y[3] Y[3] AYC[3] YM[3] AYT[3] AY[3] BIST1B BIST2 CK1B CK2 VDDHD VDDI 
+ VSSI S1BSVTSWSO8000Y24_ABUF_WOBIST
XIDEC_CKD CKPDCLK CLK_DR CKD EN_DCLK ENC WEB3B VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1_DCLK
XCKBUF CK1B CK2 CKP CLK VDDHD VDDI VSSI S1BSVTSWSO8000Y24_CKBUF_M8_DR
XABUF_PDEC_X2 AX[6] AX[7] BIST1B BIST2 CK1B CK2 X[6] X[7] XM[6] XM[7] XC[0] 
+ XC[1] XC[2] XC[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_ABUF_DECB2_WOBIST
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 EN ENC EN_D EN_DCLK RSC VDDHD VDDI VSSI 
+ S1BSVTSWSO8000Y24_ENBUFB_M8_WOBIST
XI27 AYC[3] VSSI VSSI VDDHD VDDI AYC1B[3] S1BSVTSWSO8000Y24_INV_BULK FN=3 WN=0.2U LN=0.03U 
+ MULTI=1 FP=3 WP=0.3U LP=0.03U
XI303 WEB3B VSSI VSSI VDDHD VDDI WEB4 S1BSVTSWSO8000Y24_INV_BULK FN=3 WN=0.2U LN=0.03U MULTI=1 
+ FP=3 WP=0.3U LP=0.03U
XABUF_PDEC_Y AY[0] AY[1] AY[2] BIST1B BIST2 CK1B CK2 Y[0] Y[1] Y[2] YM[0] 
+ YM[1] YM[2] XY[0] XY[1] XY[2] XY[3] XY[4] XY[5] XY[6] XY[7] VDDHD VDDI VSSI 
+ S1BSVTSWSO8000Y24_ABUF_DECB4_WOBIST
XABUF_PDEC_X0 AX[0] AX[1] AX[2] BIST1B BIST2 CK1B CK2 X[0] X[1] X[2] XM[0] 
+ XM[1] XM[2] XA[0] XA[1] XA[2] XA[3] XA[4] XA[5] XA[6] XA[7] VDDHD VDDI VSSI 
+ S1BSVTSWSO8000Y24_ABUF_DECB4_WOBIST
XABUF_PDEC_X1 AX[3] AX[4] AX[5] BIST1B BIST2 CK1B CK2 X[3] X[4] X[5] XM[3] 
+ XM[4] XM[5] XB[0] XB[1] XB[2] XB[3] XB[4] XB[5] XB[6] XB[7] VDDHD VDDI VSSI 
+ S1BSVTSWSO8000Y24_ABUF_DECB4_WOBIST
XABUF_PDEC_X3 AX[8] AX[9] AX[10] BIST1B BIST2 CK1B CK2 X[8] X[9] X[10] XM[8] 
+ XM[9] XM[10] Z[0] Z[1] Z[2] Z[3] Z[4] Z[5] Z[6] Z[7] VDDHD VDDI VSSI 
+ S1BSVTSWSO8000Y24_ABUF_DECB4_WOBIST
XIDEC_X3[0] CKP CLK_DR DEC_X3[0] EN ENC Z[0] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1_BS_SEG
XIDEC_X3[1] CKP CLK_DR DEC_X3[1] EN ENC Z[1] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1_BS_SEG
XIDEC_X3[2] CKP CLK_DR DEC_X3[2] EN ENC Z[2] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1_BS_SEG
XIDEC_X3[3] CKP CLK_DR DEC_X3[3] EN ENC Z[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1_BS_SEG
XIDEC_X3[4] CKP CLK_DR DEC_X3[4] EN ENC Z[4] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1_BS_SEG
XIDEC_X3[5] CKP CLK_DR DEC_X3[5] EN ENC Z[5] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1_BS_SEG
XIDEC_X3[6] CKP CLK_DR DEC_X3[6] EN ENC Z[6] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1_BS_SEG
XIDEC_X3[7] CKP CLK_DR DEC_X3[7] EN ENC Z[7] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_DECB1_BS_SEG
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    VHILO_V2_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_VHILO_V2_M8 VDDI VHI VLO VSSI
*.PININFO VHI:O VLO:O VDDI:B VSSI:B
MN3 VSSI Z2 Z1 VSSI nch_mac L=30N W=360N M=1
MN0 VSSI Z1 Z1 VSSI nch_mac L=30N W=360N M=1
MN1 VSSI Z2 VLO VSSI nch_mac L=30N W=1U M=3
MP7 Z2 Z1 VDDI VDDI pch_mac L=30N W=360N M=1
MP2 VHI Z1 VDDI VDDI pch_mac L=30N W=0.75U M=4
MP0 Z2 Z2 VDDI VDDI pch_mac L=30N W=360N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    CKG
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_CKG CKP CLK EN RSC RSTCK SLP_Q TM VDDHD VDDI VSSI
*.PININFO CLK:I EN:I RSTCK:I SLP_Q:I TM:I CKP:O RSC:O VDDHD:B VDDI:B VSSI:B
XINV0_MIXV_SLH SLP_Q Z17 VSSI VSSI VDDHD VDDI RSC S1BSVTSWSO8000Y24_NOR_BULK FN1=2 WN1=0.375U 
+ LN1=0.03U FN2=2 WN2=0.375U LN2=0.03U FP2=3 WP2=0.54U LP2=0.03U MULTI=1 FP1=2 
+ WP1=0.57U LP1=0.03U
XNAND0_MIXV_SLH TM CLK VSSI VSSI VDDHD VDDI Z15 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.27U 
+ LN1=0.03U FN2=1 WN2=0.27U LN2=0.03U FP2=1 WP2=0.2U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.2U LP1=0.03U
XNAND3_MIXV_SLH Z14 Z16 VSSI VSSI VDDHD VDDI Z17 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.32U 
+ LN1=0.03U FN2=1 WN2=0.32U LN2=0.03U FP2=1 WP2=0.27U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.27U LP1=0.03U
XNAND5_MIXV_SSH CKP RSC VSSI VSSI VDDHD VDDI Z19 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.27U 
+ LN1=0.03U FN2=1 WN2=0.27U LN2=0.03U FP2=1 WP2=0.5U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.375U LP1=0.03U
XNAND2_MIXV_SLH Z17 CLK VSSI VSSI VDDHD VDDI Z14 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.2U 
+ LN1=0.03U FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.2U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.2U LP1=0.03U
XNAND4_MIXV_SSH Z19 CKPC VSSI VSSI VDDHD VDDI CKP S1BSVTSWSO8000Y24_NAND_BULK FN1=3 WN1=0.67U 
+ LN1=0.03U FN2=3 WN2=0.67U LN2=0.03U FP2=2 WP2=1.1U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.2U LP1=0.03U
XNAND1_MIXV_SLH Z15 CKP RSTCK VSSI VSSI VDDHD VDDI Z16 S1BSVTSWSO8000Y24_NAND3_BULK FN1=1 
+ WN1=0.27U LN1=0.03U FN2=2 WN2=0.27U LN2=0.03U FN3=1 WN3=0.27U LN3=0.03U 
+ FP3=1 WP3=0.2U LP3=0.03U FP2=2 WP2=0.2U LP2=0.03U MULTI=1 FP1=1 WP1=0.2U 
+ LP1=0.03U
XNAND12_MIXV_SSH RSC EN CLK VSSI VSSI VDDHD VDDI CKPC S1BSVTSWSO8000Y24_NAND3_BULK FN1=1 
+ WN1=0.54U LN1=0.03U FN2=1 WN2=1.125U LN2=0.03U FN3=1 WN3=1.125U LN3=0.03U 
+ FP3=1 WP3=0.54U LP3=0.03U FP2=1 WP2=0.54U LP2=0.03U MULTI=1 FP1=1 WP1=0.75U 
+ LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    AWTD_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_AWTD_M8 AWT AWT2 VDDHD VDDI VSSI
*.PININFO AWT:I AWT2:O VDDHD:B VDDI:B VSSI:B
XINV1 AWT VSSI VSSI VDDHD VDDI NET20 S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=750N LN=0.03U MULTI=1 
+ FP=3 WP=760N LP=0.03U
MM0 AWT2 NET20 VDDHD VDDI pch_mac L=30N W=0.62U M=6
MM1 AWT2 NET20 VDDHD VDDI pch_mac L=30N W=0.76U M=7
MM2 AWT2 NET20 VSSI VSSI nch_mac L=30N W=0.75U M=8
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    RESETD_TSEL_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_RESETD_TSEL_M8 CKP V[0] V[1] VDDHD VDDI VSSI TD_01_11 TD_10
*.PININFO CKP:I V[0]:I V[1]:I TD_01_11:O TD_10:O VDDHD:B VDDI:B VSSI:B
MM10_MIXV_SSH NET75 Z4 VSSI VSSI nch_mac L=30N W=120N M=1
MM9_MIXV_SSH Z5 Z4 NET75 VSSI nch_mac L=30N W=120N M=1
MM3_MIXV_SSH NET59 Z3 VSSI VSSI nch_mac L=30N W=120N M=1
MM2_MIXV_SSH Z4 Z3 NET59 VSSI nch_mac L=30N W=120N M=1
MM22_MIXV_SSH NET43 CKP VSSI VSSI nch_mac L=30N W=120N M=1
MM16_MIXV_SSH Z3 CKP NET43 VSSI nch_mac L=30N W=120N M=1
MM8_MIXV_SSH NET83 Z4 VDDHD VDDI pch_mac L=30N W=150N M=1
MM7_MIXV_SSH Z5 Z4 NET78 VDDI pch_mac L=30N W=150N M=1
MM6_MIXV_SSH NET78 Z4 NET83 VDDI pch_mac L=30N W=150N M=1
MM5_MIXV_SSH NET84 Z3 VDDHD VDDI pch_mac L=30N W=150N M=1
MM0_MIXV_SSH Z4 Z3 NET62 VDDI pch_mac L=30N W=150N M=1
MM1_MIXV_SSH NET62 Z3 NET84 VDDI pch_mac L=30N W=150N M=1
MM4_MIXV_SSH NET85 CKP VDDHD VDDI pch_mac L=30N W=150N M=1
MM31_MIXV_SSH NET46 CKP NET85 VDDI pch_mac L=30N W=150N M=1
MM30_MIXV_SSH Z3 CKP NET46 VDDI pch_mac L=30N W=150N M=1
XND5_MIXV_SSH Z5 V[1] VSSI VSSI VDDHD VDDI TD_10 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.15U 
+ LN1=0.03U FN2=1 WN2=0.15U LN2=0.03U FP2=1 WP2=0.15U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.15U LP1=0.03U
XND1_MIXV_SSH Z0 V[0] VSSI VSSI VDDHD VDDI TD_01_11 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 
+ WN1=0.12U LN1=0.03U FN2=1 WN2=0.12U LN2=0.03U FP2=1 WP2=0.12U LP2=0.03U 
+ MULTI=1 FP1=1 WP1=0.12U LP1=0.03U
XND0_MIXV_SSH CKP TD_10 VSSI VSSI VDDHD VDDI Z0 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.12U 
+ LN1=0.03U FN2=1 WN2=0.12U LN2=0.03U FP2=1 WP2=0.12U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.12U LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    RESETD_M8_V2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_RESETD_M8_V2 BLTRKWLDRV CK2 CKP CKPD CKPDCLK IOSAEB RSTCK TK TRKBL 
+ VDDHD VDDI VSSI WEBXL WLP_SAE WLP_SAE_TK PTSEL RV[0] RV[1] WV[0] WV[1] WV[2]
*.PININFO CK2:I CKP:I WEBXL:I PTSEL:I RV[0]:I RV[1]:I WV[0]:I WV[1]:I WV[2]:I 
*.PININFO BLTRKWLDRV:O CKPD:O CKPDCLK:O IOSAEB:O RSTCK:O WLP_SAE:O TK:B 
*.PININFO TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XI622 CKP RV[0] RV[1] VDDHD VDDI VSSI RTD_01_11 RTD_10 S1BSVTSWSO8000Y24_RESETD_TSEL_M8
XI591_MIXV_SSH TRKBL2B VSSI VSSI VDDHD VDDI TRKBL3B S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=300N 
+ LN=30N MULTI=1 FP=2 WP=200N LP=30N
XI53_MIXV_SSH TRKBL VSSI VSSI VDDHD VDDI TRKBL1B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=300N 
+ LN=30N MULTI=1 FP=1 WP=300N LP=30N
XI001_MIXV_SSH NET0243 VSSI VSSI VDDHD VDDI NET0237 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=150N 
+ LN=30N MULTI=1 FP=1 WP=150N LP=30N
XI534 NET342 VSSI VSSI VDDHD VDDI NET327 S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.2U LN=0.03U 
+ MULTI=1 FP=2 WP=0.3U LP=0.03U
XI537 NET0440 VSSI VSSI VDDHD VDDI BLTRKWLDRV S1BSVTSWSO8000Y24_INV_BULK FN=8 WN=325N LN=35N 
+ MULTI=1 FP=8 WP=660N LP=35N
XINV1 TRKBL2 VSSI VSSI VDDHD VDDI Z0 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.1U LN=0.03U MULTI=1 
+ FP=1 WP=0.15U LP=0.03U
XINV0 CKP VSSI VSSI VDDHD VDDI Z6 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.12U LP=0.03U
XI533 NET327 VSSI VSSI VDDHD VDDI NET299 S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.75U LN=0.03U 
+ MULTI=1 FP=2 WP=1.125U LP=0.03U
XI507 WLP_SAE VSSI VSSI VDDHD VDDI TRKBL4 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XI566 WLP_SAE_TK VSSI VSSI VDDHD VDDI WLP_SAE_TK1B S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.6U 
+ LN=0.03U MULTI=1 FP=2 WP=0.3U LP=0.03U
XINV8 Z10 VSSI VSSI VDDHD VDDI CKPDCLK S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.75U LN=0.03U 
+ MULTI=1 FP=1 WP=1.125U LP=0.03U
XINV7 CKPD VSSI VSSI VDDHD VDDI Z10 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U LN=0.03U MULTI=1 
+ FP=1 WP=0.3U LP=0.03U
XINV6 Z8 VSSI VSSI VDDHD VDDI CKPD S1BSVTSWSO8000Y24_INV_BULK FN=4 WN=0.75U LN=0.03U MULTI=1 
+ FP=4 WP=1.125U LP=0.03U
XINV5 CKP VSSI VSSI VDDHD VDDI Z8 S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=300N LN=0.03U MULTI=1 
+ FP=2 WP=400N LP=0.03U
XI532 NET299 VSSI VSSI VDDHD VDDI IOSAEB S1BSVTSWSO8000Y24_INV_BULK FN=5 WN=0.75U LN=0.03U 
+ MULTI=1 FP=6 WP=1.195U LP=0.03U
XI598 D6 VSSI VSSI VDDHD VDDI D7 S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.15U LN=0.03U MULTI=1 
+ FP=2 WP=0.3U LP=0.03U
XI000_MIXV_SSH CKP VSSI VSSI VDDHD VDDI NET0243 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=150N LN=30N 
+ MULTI=1 FP=1 WP=150N LP=30N
XI618_MIXV_SSH TRKBL1B VSSI VSSI VDDHD VDDI TRKBL2B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=300N 
+ LN=30N MULTI=1 FP=2 WP=200N LP=30N
MM18D_MIXV_SSH NET0194 D4 VDDHD VDDI pch_mac L=30N W=120N M=1
MM15D_MIXV_SSH NET0197 D3 VDDHD VDDI pch_mac L=30N W=120N M=1
MM14D_MIXV_SSH D4 D3 NET0197 VDDI pch_mac L=30N W=120N M=1
MM11D_MIXV_SSH D3 D2 NET0199 VDDI pch_mac L=30N W=120N M=1
MM10D_MIXV_SSH NET0199 D2 VDDHD VDDI pch_mac L=30N W=120N M=1
MM7D_MIXV_SSH NET0200 D1 VDDHD VDDI pch_mac L=30N W=120N M=1
MM6D_MIXV_SSH D2 D1 NET0200 VDDI pch_mac L=30N W=120N M=1
MM3D_MIXV_SSH NET0203 WEBXL VDDHD VDDI pch_mac L=30N W=120N M=1
MM2D_MIXV_SSH D1 WEBXL NET0203 VDDI pch_mac L=30N W=120N M=1
MM25_MIXV_SSH NET0454 Z4 VDDHD VDDI pch_mac L=30N W=120N M=1
MM24_MIXV_SSH Z5 NET0454 NET0396 VDDI pch_mac L=30N W=120N M=1
MM23_MIXV_SSH NET0396 NET0454 VDDHD VDDI pch_mac L=30N W=120N M=1
MM19D_MIXV_SSH D5 D4 NET0194 VDDI pch_mac L=30N W=120N M=1
MM7_MIXV_SSH NET0494 NET0415 VDDHD VDDI pch_mac L=30N W=120N M=1
MM16_MIXV_SSH NET0474 Z3 VDDHD VDDI pch_mac L=30N W=120N M=1
MM20_MIXV_SSH NET0408 NET0474 VDDHD VDDI pch_mac L=30N W=120N M=1
MM23D_MIXV_SSH D6 D5 NET0192 VDDI pch_mac L=30N W=120N M=1
MM22D_MIXV_SSH NET0192 D5 VDDHD VDDI pch_mac L=30N W=120N M=1
MM5_MIXV_SSH NET0415 WLP_SAE NET0401 VDDI pch_mac L=30N W=120N M=1
MP16 WLP_SAE TRKBL2 VDDHD VDDI pch_mac L=30N W=1.2U M=5
MP161 WLP_SAE TRKBL2 VDDHD VDDI pch_mac L=30N W=1.125U M=6
MM12_MIXV_SSH Z3 NET0494 NET0420 VDDI pch_mac L=30N W=120N M=1
MM19_MIXV_SSH Z4 NET0474 NET0408 VDDI pch_mac L=30N W=120N M=1
MM11_MIXV_SSH NET0420 NET0494 VDDHD VDDI pch_mac L=30N W=120N M=1
MM3_MIXV_SSH NET0401 WLP_SAE VDDHD VDDI pch_mac L=30N W=120N M=1
MM17D_MIXV_SSH NET0195 D4 VSSI VSSI nch_mac L=30N W=120N M=1
MM16D_MIXV_SSH D5 D4 NET0195 VSSI nch_mac L=30N W=120N M=1
MM13D_MIXV_SSH D4 D3 NET0196 VSSI nch_mac L=30N W=120N M=1
MM12D_MIXV_SSH NET0196 D3 VSSI VSSI nch_mac L=30N W=120N M=1
MM9D_MIXV_SSH D3 D2 NET0198 VSSI nch_mac L=30N W=120N M=1
MM8D_MIXV_SSH NET0198 D2 VSSI VSSI nch_mac L=30N W=120N M=1
MM5D_MIXV_SSH NET0201 D1 VSSI VSSI nch_mac L=30N W=120N M=1
MM4D_MIXV_SSH D2 D1 NET0201 VSSI nch_mac L=30N W=120N M=1
MM1D_MIXV_SSH D1 WEBXL NET0202 VSSI nch_mac L=30N W=120N M=1
MM30_MIXV_SSH NET0450 Z4 VSSI VSSI nch_mac L=30N W=120N M=1
MM29_MIXV_SSH NET0454 Z4 NET0450 VSSI nch_mac L=30N W=120N M=1
MM28_MIXV_SSH Z5 NET0454 VSSI VSSI nch_mac L=30N W=120N M=1
MM21_MIXV_SSH Z4 NET0474 VSSI VSSI nch_mac L=30N W=120N M=1
MM17_MIXV_SSH NET0478 Z3 VSSI VSSI nch_mac L=30N W=120N M=1
MM14_MIXV_SSH Z3 NET0494 VSSI VSSI nch_mac L=30N W=120N M=1
MM9_MIXV_SSH NET0494 NET0415 NET0490 VSSI nch_mac L=30N W=120N M=1
MM6_MIXV_SSH NET0415 WLP_SAE VSSI VSSI nch_mac L=30N W=120N M=1
MM21D_MIXV_SSH D6 D5 NET0193 VSSI nch_mac L=30N W=120N M=1
MM20D_MIXV_SSH NET0193 D5 VSSI VSSI nch_mac L=30N W=120N M=1
MN7 WLP_SAE TRKBL2 VSSI VSSI nch_mac L=30N W=0.375U M=12
MM18_MIXV_SSH NET0474 Z3 NET0478 VSSI nch_mac L=30N W=120N M=1
MM10_MIXV_SSH NET0490 NET0415 VSSI VSSI nch_mac L=30N W=120N M=1
MM0D_MIXV_SSH NET0202 WEBXL VSSI VSSI nch_mac L=30N W=120N M=1
XNAND3 CKP RTD_10 RTD_01_11 VSSI VSSI VDDHD VDDI NET0440 S1BSVTSWSO8000Y24_NAND3_BULK FN1=2 
+ WN1=1.145U LN1=30N FN2=2 WN2=1.145U LN2=30N FN3=2 WN3=1.145U LN3=30N FP3=2 
+ WP3=400N LP3=30N FP2=2 WP2=400N LP2=30N MULTI=1 FP1=2 WP1=400N LP1=30N
XI521 TRKBL2 WLP_SAE_TK1B Z5 VSSI VSSI VDDHD VDDI NET342 S1BSVTSWSO8000Y24_NAND3_BULK FN1=1 
+ WN1=0.4U LN1=0.03U FN2=1 WN2=0.4U LN2=0.03U FN3=1 WN3=0.4U LN3=0.03U FP3=1 
+ WP3=0.3U LP3=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 WP1=0.3U LP1=0.03U
XTSEL_WT TRKBL1B TK VDDHD VDDI VSSI NET0313 WV[0] WV[1] S1BSVTSWSO8000Y24_RESETD_TSEL_WT
XI12_MIXV_SSH RSTCKB Z8 VSSI VSSI VDDHD VDDI RSTCK S1BSVTSWSO8000Y24_NOR_BULK FN1=1 WN1=0.2U 
+ LN1=0.03U FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.6U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.6U LP1=0.03U
XI574_MIXV_SSH NET0313 TRKBL1B VSSI VSSI VDDHD VDDI RSTCKB S1BSVTSWSO8000Y24_NAND_BULK FN1=1 
+ WN1=0.45U LN1=30N FN2=1 WN2=0.45U LN2=30N FP2=1 WP2=400N LP2=30N MULTI=1 
+ FP1=1 WP1=400N LP1=30N
XI587 D7 TRKBL3B VSSI VSSI VDDHD VDDI TRKBL2 S1BSVTSWSO8000Y24_NAND_BULK FN1=4 WN1=1U 
+ LN1=0.03U FN2=4 WN2=1U LN2=0.03U FP2=2 WP2=1U LP2=0.03U MULTI=1 FP1=2 WP1=1U 
+ LP1=0.03U
XNAND0 Z6 Z6 VSSI VSSI VDDHD VDDI Z7 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.2U LN1=0.03U 
+ FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 WP1=0.3U 
+ LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    COTH_M8_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_COTH_M8_WOBIST AWT AWT2 BLTRKWLDRV CK2 CKP CKPD CKPDCLK CLK DSLP 
+ DSLP_BUF EN PTSEL RSC RTSEL[0] RTSEL[1] SD SD_BUF SLP SLP_BUF SLP_Q TK TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WEB3B WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2]
*.PININFO AWT:I CK2:I CLK:I DSLP:I EN:I PTSEL:I RTSEL[0]:I RTSEL[1]:I SD:I 
*.PININFO SLP:I SLP_Q:I TM:I WEB3B:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I AWT2:O 
*.PININFO BLTRKWLDRV:O CKP:O CKPD:O CKPDCLK:O DSLP_BUF:O RSC:O SD_BUF:O 
*.PININFO SLP_BUF:O VHI:O VLO:O WLP_SAE:O WLP_SAEB:O TK:B TRKBL:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WLP_SAE_TK:B
XVHILO VDDI VHI VLO VSSI S1BSVTSWSO8000Y24_VHILO_V2_M8
XPMCTRL CKP DSLP DSLP_BUF SD SD_BUF SLP SLP_BUF VDDI VSSI S1BSVTSWSO8000Y24_PMCTRL
XCKG CKP CLK EN RSC RSTCK SLP_Q TM VDDHD VDDI VSSI S1BSVTSWSO8000Y24_CKG
XAWTD AWT AWT2 VDDHD VDDI VSSI S1BSVTSWSO8000Y24_AWTD_M8
XRESETD BLTRKWLDRV CK2 CKP CKPD CKPDCLK WLP_SAEB RSTCK TK TRKBL VDDHD VDDI 
+ VSSI WEB3B WLP_SAE WLP_SAE_TK PTSEL RTSEL[0] RTSEL[1] WTSEL[0] WTSEL[1] 
+ WTSEL[2] S1BSVTSWSO8000Y24_RESETD_M8_V2
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    CNT_CORE_M16_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_CNT_CORE_M16_WOBIST AWT AWT2 BLTRKWLDRV CEB CEBM CKD CLK CLK_DR 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP 
+ DSLP_BUF PTSEL RE REDEN REDENB RTSEL[0] RTSEL[1] SD SD_BUF SLP SLP_BUF SLP_Q 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] 
+ X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] 
+ Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I CEB:I CEBM:I CLK:I CLK_DR:I DSLP:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I SD:I SLP:I SLP_Q:I TM:I WEB:I WEBM:I 
*.PININFO WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I 
*.PININFO X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I 
*.PININFO XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O DSLP_BUF:O RE:O SD_BUF:O SLP_BUF:O VHI:O VLO:O WE:O 
*.PININFO WLP_SAE:O WLP_SAEB:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B 
*.PININFO VSSI:B WLP_SAE_TK:B
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK2 CKD CKP CKPD CKPDCLK CLK CLK_DR DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] 
+ DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] 
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN RE REDEN 
+ REDENB RSC VDDHD VDDI VSSI WE WEB WEB3B WEBM X[0] X[1] X[2] X[3] X[4] X[5] 
+ X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1BSVTSWSO8000Y24_CDEC_M8_WOBIST
XCOTHERS AWT AWT2 BLTRKWLDRV CKP CKP CKPD CKPDCLK CLK DSLP DSLP_BUF EN PTSEL 
+ RSC RTSEL[0] RTSEL[1] SD SD_BUF SLP SLP_BUF SLP_Q TK TM TRKBL VDDHD VDDI VHI 
+ VLO VSSI WEB3B WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1BSVTSWSO8000Y24_COTH_M8_WOBIST
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    CNT_M16_IOX2_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_CNT_M16_IOX2_WOBIST AWT AWT2 BLTRKWLDRV BWEBM_L BWEBM_R BWEB_L BWEB_R 
+ CEB CEBM CKD CLK CLK_DR DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DM_L DM_R DSLP DSLP_BUF D_L D_R GBLB_L GBLB_R GBL_L GBL_R 
+ GWB_L GWB_R GW_L GW_R PTSEL Q_L Q_R RE REDEN REDENB RTSEL[0] RTSEL[1] SD 
+ SD_BUF SLP SLP_BUF SLP_LBACK SLP_LCTRL SLP_Q SLP_RBACK TK TM TRKBL VDDF 
+ VDDFHD VDDHD VDDI VHI VLO VSSI WE WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] 
+ X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] 
+ Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BWEBM_L:I BWEBM_R:I BWEB_L:I BWEB_R:I CEB:I CEBM:I CLK:I 
*.PININFO CLK_DR:I DM_L:I DM_R:I DSLP:I D_L:I D_R:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I SD:I SLP:I SLP_LBACK:I SLP_RBACK:I TM:I WEB:I 
*.PININFO WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I 
*.PININFO X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I 
*.PININFO XM[10]:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I 
*.PININFO GWB_L:O GWB_R:O GW_L:O GW_R:O Q_L:O Q_R:O SLP_LCTRL:O SLP_Q:O AWT2:B 
*.PININFO BLTRKWLDRV:B CKD:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DSLP_BUF:B GBLB_L:B GBLB_R:B GBL_L:B GBL_R:B RE:B 
*.PININFO SD_BUF:B SLP_BUF:B TK:B TRKBL:B VDDF:B VDDFHD:B VDDHD:B VDDI:B VHI:B 
*.PININFO VLO:B VSSI:B WE:B WLP_SAE:B WLP_SAEB:B WLP_SAE_TK:B YL[0]:B YL[1]:B
MM4 VDDHD SLP_BUF VDDI VDDI pch_mac L=35.0N W=1U M=5
MM2 VDDHD SLP_BUF VDDI VDDI pch_mac L=35.0N W=0.75U M=16
MM1 VDDHD SLP_BUF VDDI VDDI pch_mac L=35.0N W=0.4U M=8
MM0 VDDHD SLP_BUF VDDI VDDI pch_mac L=35.0N W=1U M=70
XI14 SLP_RBACK SLP_LBACK VSSI VSSI VDDI VDDI NET158 S1BSVTSWSO8000Y24_NOR_BULK FN1=1 WN1=0.3U 
+ LN1=0.035U FN2=1 WN2=0.3U LN2=0.035U FP2=1 WP2=0.6U LP2=0.035U MULTI=1 FP1=1 
+ WP1=0.6U LP1=0.035U
XI17 NET158 VSSI VSSI VDDI VDDI SLP_LCTRL S1BSVTSWSO8000Y24_INV_BULK FN=6 WN=0.3U LN=0.035U 
+ MULTI=1 FP=6 WP=0.6U LP=0.035U
XI15 NET158 VSSI VSSI VDDI VDDI SLP_Q S1BSVTSWSO8000Y24_INV_BULK FN=4 WN=0.3U LN=0.035U 
+ MULTI=1 FP=4 WP=0.6U LP=0.035U
MM9[0] DEC_X0[0] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM9[1] DEC_X0[1] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM9[2] DEC_X0[2] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM9[3] DEC_X0[3] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM9[4] DEC_X0[4] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM9[5] DEC_X0[5] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM9[6] DEC_X0[6] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM9[7] DEC_X0[7] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM5[0] DEC_X1[0] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM5[1] DEC_X1[1] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM5[2] DEC_X1[2] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM5[3] DEC_X1[3] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM5[4] DEC_X1[4] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM5[5] DEC_X1[5] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM5[6] DEC_X1[6] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
MM5[7] DEC_X1[7] SLP_Q VSSI VSSI nch_mac L=30N W=140N M=1
XIO_R AWT2 BWEB_R BWEBM_R CKD D_R DM_R GBL_R GBLB_R GW_R GWB_R Q_R SLP_Q VDDF 
+ VDDFHD VDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_WOBIST
XIO_L AWT2 BWEB_L BWEBM_L CKD D_L DM_L GBL_L GBLB_L GW_L GWB_L Q_L SLP_Q VDDF 
+ VDDFHD VDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_WOBIST
XCNT AWT AWT2 BLTRKWLDRV CEB CEBM CKD CLK CLK_DR DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] VLO DSLP_BUF PTSEL RE REDEN REDENB 
+ RTSEL[0] RTSEL[1] SD SD_BUF SLP SLP_BUF SLP_Q TK TM TRKBL VDDHD VDDI VHI VLO 
+ VSSI WE WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] 
+ XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] 
+ YM[0] YM[1] YM[2] YM[3] S1BSVTSWSO8000Y24_CNT_CORE_M16_WOBIST
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    XDRV_STRAP
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_XDRV_STRAP VDDHD VDDI VSSI WLPY WLPYB
*.PININFO WLPY:I VDDHD:B VDDI:B VSSI:B WLPYB:B
MN1 WLPYB WLPY VSSI VSSI nch_mac L=30N W=0.8U M=10
MP0 WLPYB WLPY VDDHD VDDI pch_mac L=30N W=0.72U M=5
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    LIO_HEADER_N1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_LIO_HEADER_N1 LIOPD PDI PDO PDO_BACK VDDAI VDDI VSSI
*.PININFO LIOPD:I PDI:I PDO_BACK:I PDO:O VDDAI:B VDDI:B VSSI:B
XI0 NET16 VSSI VSSI VDDI VDDI PDO S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.035U MULTI=1 
+ FP=1 WP=0.12U LP=0.035U
XI1 PDI LIOPD VSSI VSSI VDDI VDDI NET16 S1BSVTSWSO8000Y24_NOR_BULK FN1=1 WN1=0.12U LN1=0.035U 
+ FN2=1 WN2=0.12U LN2=0.035U FP2=1 WP2=0.12U LP2=0.035U MULTI=1 FP1=1 
+ WP1=0.12U LP1=0.035U
MM0 VDDAI PDO_BACK VDDI VDDI pch_mac L=35.0N W=0.95U M=5
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    PRECHARGE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_PRECHARGE BL BLB BLEQB VDDAI VDDI
*.PININFO BLEQB:I BL:B BLB:B VDDAI:B VDDI:B
MP0_MIXV_SLH VDDAI BLEQB BL VDDI pch_mac L=30N W=0.44U M=3
MP5_MIXV_SLH BL BLEQB BLB VDDI pch_mac L=30N W=440N M=1
MP17_MIXV_SLH BLB BLEQB VDDAI VDDI pch_mac L=30N W=0.44U M=3
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    TKBL_BCELL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_TKBL_BCELL BLB BL_TK G_FLOAT VDDAI VDDI VSSI WL WL_TK TIEH
*.PININFO WL:I WL_TK:I BLB:B BL_TK:B G_FLOAT:B VDDAI:B VDDI:B VSSI:B TIEH:B
MPCHPU1 TIEH BL_TK_IN VDDAI VDDI pchpu_sr L=35N W=40N M=1
MPCHPU0 VDDAI TIEH BL_TK_IN VDDI pchpu_sr L=35N W=40N M=1
MNCHPD1 TIEH BL_TK_IN G_FLOAT VSSI nchpd_sr L=35N W=95N M=1
MNCHPD0 VSSI TIEH BL_TK_IN VSSI nchpd_sr L=35N W=95N M=1
MNCHPG1 TIEH WL BLB VSSI nchpg_sr L=35N W=65N M=1
MNCHPG0 BL_TK WL_TK BL_TK_IN VSSI nchpg_sr L=35N W=65N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    TRKNOR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_TRKNOR BLB BLB_EDGE BL_EDGE BL_TK G_FLOAT VDDAI VDDI VSSI WL WL_TK TIEH
*.PININFO WL:I WL_TK:I TIEH:I BLB:B BLB_EDGE:B BL_EDGE:B BL_TK:B G_FLOAT:B 
*.PININFO VDDAI:B VDDI:B VSSI:B
XTKBL_BCELL BLB BL_TK G_FLOAT VDDAI VDDI VSSI WL WL_TK TIEH S1BSVTSWSO8000Y24_TKBL_BCELL
XTKBL_BCELL_RIGHT BLB_EDGE BL_EDGE G_FLOAT VDDAI VDDI VSSI WL WL_TK TIEH 
+ S1BSVTSWSO8000Y24_TKBL_EDGE
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    TRKNORX2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_TRKNORX2 BL_TK VDDAI VDDI VSSI WL[0] WL[1] WL_TK FLOAT1 FLOAT2 FLOAT3 
+ FLOAT4 FLOAT5 TIEH
*.PININFO WL[0]:I WL[1]:I WL_TK:I TIEH:I BL_TK:B VDDAI:B VDDI:B VSSI:B 
*.PININFO FLOAT1:B FLOAT2:B FLOAT3:B FLOAT4:B FLOAT5:B
XTRKNOR_1 FLOAT2 FLOAT4 FLOAT1 BL_TK G_FLOAT VDDAI VDDI VSSI WL[1] WL_TK TIEH 
+ S1BSVTSWSO8000Y24_TRKNOR
XTRKNOR_0 FLOAT3 FLOAT5 FLOAT1 BL_TK G_FLOAT VDDAI VDDI VSSI WL[0] WL_TK TIEH 
+ S1BSVTSWSO8000Y24_TRKNOR
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    MCB_TKWL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_MCB_TKWL BL BLB VDDAI VDDI VSSI WL
*.PININFO BL:B BLB:B VDDAI:B VDDI:B VSSI:B WL:B
MPCHPU1 VSSI BL_IN P_FLOAT VDDI pchpu_sr L=35N W=40N M=1
MPCHPU0 VDDAI VSSI BL_IN VDDI pchpu_sr L=35N W=40N M=1
MNCHPD1 VSSI BL_IN VSSI VSSI nchpd_sr L=35N W=95N M=1
MNCHPD0 VSSI VSSI BL_IN VSSI nchpd_sr L=35N W=95N M=1
MNCHPG1 BLB WL VSSI VSSI nchpg_sr L=35N W=65N M=1
MNCHPG0 BL_IN WL BL VSSI nchpg_sr L=35N W=65N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    MCB_TKWL_ISO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_MCB_TKWL_ISO BL BLB VDDAI VDDI VSSI WLL WLR
*.PININFO BL:B BLB:B VDDAI:B VDDI:B VSSI:B WLL:B WLR:B
MNCHPG1 BLB WLR VSSI VSSI nchpg_sr L=35N W=65N M=1
MNCHPG0 NET060 WLL BL VSSI nchpg_sr L=35N W=65N M=1
MNCHPD1 VSSI NET060 VSSI VSSI nchpd_sr L=35N W=95N M=1
MNCHPD0 VSSI VSSI NET060 VSSI nchpd_sr L=35N W=95N M=1
MPCHPU1 VSSI NET060 P_FLOAT VDDI pchpu_sr L=35N W=40N M=1
MPCHPU0 VDDAI VSSI NET060 VDDI pchpu_sr L=35N W=40N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    TKWL_2X2_ISO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_TKWL_2X2_ISO VDDAI VDDI VSSI WL_TK_L[0] WL_TK_L[1] WL_TK_R[0] 
+ WL_TK_R[1]
*.PININFO WL_TK_L[0]:I WL_TK_L[1]:I WL_TK_R[0]:I WL_TK_R[1]:I VDDAI:B VDDI:B 
*.PININFO VSSI:B
XI25 NET294 NET278 VDDAI VDDI VSSI WL_TK_R[0] WL_TK_L[0] S1BSVTSWSO8000Y24_MCB_TKWL_ISO
XI22 NET279 NET278 VDDAI VDDI VSSI WL_TK_R[1] WL_TK_L[1] S1BSVTSWSO8000Y24_MCB_TKWL_ISO
XI24 NET030 NET284 VDDAI VDDI VSSI WL_TK_R[0] S1BSVTSWSO8000Y24_MCB_TKWL
XTKWL_MCB_1 NET281 NET284 VDDAI VDDI VSSI WL_TK_R[1] S1BSVTSWSO8000Y24_MCB_TKWL
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    MCB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_MCB BL BLB VDDAI VDDI VSSI WL
*.PININFO BL:B BLB:B VDDAI:B VDDI:B VSSI:B WL:B
MPCHPU1 BLB_IN BL_IN VDDAI VDDI pchpu_sr L=35N W=40N M=1
MPCHPU0 VDDAI BLB_IN BL_IN VDDI pchpu_sr L=35N W=40N M=1
MNCHPD1 BLB_IN BL_IN VSSI VSSI nchpd_sr L=35N W=95N M=1
MNCHPD0 VSSI BLB_IN BL_IN VSSI nchpd_sr L=35N W=95N M=1
MNCHPG1 BLB WL BLB_IN VSSI nchpg_sr L=35N W=65N M=1
MNCHPG0 BL_IN WL BL VSSI nchpg_sr L=35N W=65N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    MCB_2X16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_MCB_2X16 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] 
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] 
+ BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] 
+ BLB[15] GBL GBLB GW GWB VDDAI VDDI VSSI WL[0] WL[1]
*.PININFO BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B BL[6]:B BL[7]:B 
*.PININFO BL[8]:B BL[9]:B BL[10]:B BL[11]:B BL[12]:B BL[13]:B BL[14]:B 
*.PININFO BL[15]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B BLB[5]:B 
*.PININFO BLB[6]:B BLB[7]:B BLB[8]:B BLB[9]:B BLB[10]:B BLB[11]:B BLB[12]:B 
*.PININFO BLB[13]:B BLB[14]:B BLB[15]:B GBL:B GBLB:B GW:B GWB:B VDDAI:B VDDI:B 
*.PININFO VSSI:B WL[0]:B WL[1]:B
XMCB_1[0] BL[0] BLB[0] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[1] BL[1] BLB[1] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[2] BL[2] BLB[2] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[3] BL[3] BLB[3] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[4] BL[4] BLB[4] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[5] BL[5] BLB[5] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[6] BL[6] BLB[6] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[7] BL[7] BLB[7] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[8] BL[8] BLB[8] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[9] BL[9] BLB[9] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[10] BL[10] BLB[10] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[11] BL[11] BLB[11] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[12] BL[12] BLB[12] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[13] BL[13] BLB[13] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[14] BL[14] BLB[14] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_1[15] BL[15] BLB[15] VDDAI VDDI VSSI WL[1] S1BSVTSWSO8000Y24_MCB
XMCB_0[0] BL[0] BLB[0] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[1] BL[1] BLB[1] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[2] BL[2] BLB[2] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[3] BL[3] BLB[3] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[4] BL[4] BLB[4] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[5] BL[5] BLB[5] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[6] BL[6] BLB[6] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[7] BL[7] BLB[7] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[8] BL[8] BLB[8] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[9] BL[9] BLB[9] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[10] BL[10] BLB[10] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[11] BL[11] BLB[11] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[12] BL[12] BLB[12] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[13] BL[13] BLB[13] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[14] BL[14] BLB[14] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
XMCB_0[15] BL[15] BLB[15] VDDAI VDDI VSSI WL[0] S1BSVTSWSO8000Y24_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    TKBL_TRKPRE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_TKBL_TRKPRE SLP_BUF TRKBL TRKWL VDDAI VDDI VSSI ZH ZL
*.PININFO SLP_BUF:I TRKWL:I ZH:O ZL:O TRKBL:B VDDAI:B VDDI:B VSSI:B
MM7 ZH NET_021 VDDAI VDDI pch_mac L=30N W=910N M=1
MM8 NET_039 NET_039 VDDI VDDI pch_mac L=30N W=180N M=2
MM9 ZH NET_021 VDDAI VDDI pch_mac L=30N W=515N M=1
MP0_MIXV_SSH TRKBL TRKWL VDDI VDDI pch_mac L=30N W=0.9U M=2
MM10 ZH NET_021 VDDAI VDDI pch_mac L=30N W=835N M=1
MM11 ZH NET_021 VDDAI VDDI pch_mac L=30N W=740N M=1
MM4 NET_039 NET_021 VDDI VDDI pch_mac L=30N W=180N M=2
MM02 ZL NET_039 VSSI VSSI nch_mac L=30N W=0.5U M=2
MM01 ZL NET_039 VSSI VSSI nch_mac L=30N W=1U M=2
MM2 NET_021 NET_021 VSSI VSSI nch_mac L=30N W=360N M=1
MM3 NET_021 NET_039 VSSI VSSI nch_mac L=30N W=360N M=1
MM1 TRKWL SLP_BUF VSSI VSSI nch_mac L=30N W=120N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    XDRV_LA512_SHA_NMOS
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS DEC_X1 SH_NPD VSSI
*.PININFO DEC_X1:B SH_NPD:B VSSI:B
MN5 SH_NPD DEC_X1 VSSI VSSI nch_mac L=35.0N W=320N M=2
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    XDRV_STRAP_LCNT
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_XDRV_STRAP_LCNT VDDHD VDDI VSSI WLPY WLPYB
*.PININFO WLPY:I VDDHD:B VDDI:B VSSI:B WLPYB:B
MN1 WLPYB WLPY VSSI VSSI nch_mac L=30N W=2U M=4
MP0 WLPYB WLPY VDDHD VDDI pch_mac L=30N W=1.8U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    TKWL_2X2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_TKWL_2X2 VDDAI VDDI VSSI WL_DUM WL_TK
*.PININFO VDDAI:B VDDI:B VSSI:B WL_DUM:B WL_TK:B
XTKWL_MCB_1 FLOAT_BL_R_T FLOAT_BLB_R VDDAI VDDI VSSI WL_TK S1BSVTSWSO8000Y24_MCB_TKWL
XTKWL_MCB_0 FLOAT_BL_L_T FLOAT_BLB_L VDDAI VDDI VSSI WL_TK S1BSVTSWSO8000Y24_MCB_TKWL
XTKDUM_MCB_1 FLOAT_BL_R_B FLOAT_BLB_R VDDAI VDDI VSSI WL_DUM S1BSVTSWSO8000Y24_MCB_TKWL
XTKDUM_MCB_0 FLOAT_BL_L_B FLOAT_BLB_L VDDAI VDDI VSSI WL_DUM S1BSVTSWSO8000Y24_MCB_TKWL
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    DIO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_DIO A VSSI
*.PININFO A:B VSSI:B
DDIO VSSI A ndio AREA=0.02E-12 M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    XDRV_WLP_S_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_XDRV_WLP_S_M8 BLEQ BLEQB BS DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ SLP_LCTRL VDDHD VDDI VSSI WLPY[0] WLPY[1] WLPY[2] WLPY[3] WLP_SAE
*.PININFO BS:I DEC_X2[0]:I DEC_X2[1]:I DEC_X2[2]:I DEC_X2[3]:I SLP_LCTRL:I 
*.PININFO WLP_SAE:I BLEQ:O BLEQB:O WLPY[0]:O WLPY[1]:O WLPY[2]:O WLPY[3]:O 
*.PININFO VDDHD:B VDDI:B VSSI:B
XI558 WLP_SAE VSSI VSSI VDDHD VDDI D1 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.24U LP=0.03U
XI576 D3 VSSI VSSI VDDHD VDDI D4 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.24U LN=0.03U MULTI=1 
+ FP=1 WP=0.12U LP=0.03U
XI557 BLEQB VSSI VSSI VDDI VDDI BLEQ S1BSVTSWSO8000Y24_INV_BULK FN=6 WN=0.84U LN=0.03U MULTI=1 
+ FP=6 WP=0.84U LP=0.03U
XI575 D2 VSSI VSSI VDDHD VDDI D3 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.24U LP=0.03U
XI574 D1 VSSI VSSI VDDHD VDDI D2 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.24U LN=0.03U MULTI=1 
+ FP=1 WP=0.12U LP=0.03U
XI587 WLP_SAE VSSI VSSI VDDHD VDDI RD_RSTB S1BSVTSWSO8000Y24_INV_BULK FN=3 WN=0.21U LN=0.03U 
+ MULTI=1 FP=3 WP=0.4U LP=0.03U
XI577 D4 VSSI VSSI VDDHD VDDI D5 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.24U LP=0.03U
XI532 NET363 VSSI VSSI VDDHD VDDI WLPY[1] S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=1.1U LN=0.03U 
+ MULTI=1 FP=9 WP=1.1U LP=0.03U
XI531 NET371 VSSI VSSI VDDHD VDDI WLPY[3] S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=1.1U LN=0.03U 
+ MULTI=1 FP=9 WP=1.1U LP=0.03U
XI533 NET367 VSSI VSSI VDDHD VDDI WLPY[2] S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=1.1U LN=0.03U 
+ MULTI=1 FP=9 WP=1.1U LP=0.03U
XI534 MWL2[0] VSSI VSSI VDDHD VDDI WLPY[0] S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=1.1U LN=0.03U 
+ MULTI=1 FP=9 WP=1.1U LP=0.03U
XI592 NET383 VSSI VSSI VDDHD VDDI BLEQB S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.8U LN=0.03U 
+ MULTI=1 FP=4 WP=0.75U LP=0.03U
MM5 MWL2[0] RD_RSTB VDDHD VDDI pch_mac L=30N W=300N M=2
MMP4 NET371 RD_RSTB VDDHD VDDI pch_mac L=30N W=300N M=2
MM16 NET367 BS VDDHD VDDI pch_mac L=30N W=200N M=1
MM9 NET363 BS VDDHD VDDI pch_mac L=30N W=200N M=1
MM4 NET363 RD_RSTB VDDHD VDDI pch_mac L=30N W=300N M=2
MM20 MWL2[0] BS VDDHD VDDI pch_mac L=30N W=200N M=1
MM3 NET367 RD_RSTB VDDHD VDDI pch_mac L=30N W=300N M=2
MM15 NET371 DEC_X2[3] VDDHD VDDI pch_mac L=30N W=200N M=1
MM13 NET367 DEC_X2[2] VDDHD VDDI pch_mac L=30N W=200N M=1
MM12 MWL2[0] DEC_X2[0] VDDHD VDDI pch_mac L=30N W=200N M=1
MM10 NET363 DEC_X2[1] VDDHD VDDI pch_mac L=30N W=200N M=1
MM21 NET371 BS VDDHD VDDI pch_mac L=30N W=200N M=1
MM1 NET375 RD_RSTB VSSI VSSI nch_mac L=30N W=0.31U M=8
MM35 NET371 DEC_X2[3] SHARE VSSI nch_mac L=30N W=0.41U M=4
MM34 NET367 DEC_X2[2] SHARE VSSI nch_mac L=30N W=0.41U M=4
MM32 NET363 DEC_X2[1] SHARE VSSI nch_mac L=30N W=0.41U M=4
MM28 MWL2[0] DEC_X2[0] SHARE VSSI nch_mac L=30N W=0.41U M=4
MM36 BLEQB SLP_LCTRL VSSI VSSI nch_mac L=30N W=120N M=1
MM0 SHARE BS NET375 VSSI nch_mac L=30N W=0.31U M=8
XI551 D5 BS VSSI VSSI VDDHD VDDI NET383 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.8U LN1=0.03U 
+ FN2=1 WN2=0.8U LN2=0.03U FP2=1 WP2=0.4U LP2=0.03U MULTI=1 FP1=1 WP1=0.4U 
+ LP1=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    LCTRL_S_M8_SD
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_LCTRL_S_M8_SD BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ DSLP_BUF LIOPD RE RE_LIO SAEB SLP_LCTRL TK VDDHD VDDI VSSI WE WE_LIO 
+ WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] 
+ WLPY_UP[3] WLP_SAE WLP_SAE_TK YL[0] YL[1] YL_LIO[0] YL_LIO[1]
*.PININFO DSLP_BUF:I SLP_LCTRL:I BLEQ_DN:O BLEQ_UP:O DEC_Y_DN[0]:O 
*.PININFO DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O DEC_Y_DN[4]:O 
*.PININFO DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O DEC_Y_UP[0]:O 
*.PININFO DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O DEC_Y_UP[4]:O 
*.PININFO DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O LIOPD:O RE_LIO:O SAEB:O 
*.PININFO WE_LIO:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B RE:B TK:B VDDHD:B VDDI:B VSSI:B WE:B WLP_SAE:B 
*.PININFO WLP_SAE_TK:B YL[0]:B YL[1]:B
MM2 VDDHD SLP_LCTRL VDDI VDDI pch_mac L=35.0N W=1U M=142
XLCTRL_PM DSLP_BUF LIOPD SLP_LCTRL VDDI VSSI S1BSVTSWSO8000Y24_LCTRL_PM
XXDRV_WLP_DN BLEQ_DN BLEQB_DN DEC_X3[0] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] SLP_LCTRL VDDHD VDDI VSSI WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] 
+ WLPY_DN[3] WLP_SAE S1BSVTSWSO8000Y24_XDRV_WLP_S_M8
XXDRV_WLP_UP BLEQ_UP BLEQB_UP DEC_X3[1] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] SLP_LCTRL VDDHD VDDI VSSI WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] 
+ WLPY_UP[3] WLP_SAE S1BSVTSWSO8000Y24_XDRV_WLP_S_M8
XLCTRL BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] SLP_LCTRL RE RE_LIO SAEB VDDHD VDDI VSSI WE WE_LIO 
+ WLP_SAE YL[0] YL[1] YL_LIO[0] YL_LIO[1] S1BSVTSWSO8000Y24_LCTRL
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    LCTRL_S_M16_SD
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_LCTRL_S_M16_SD BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ DSLP_BUF LIOPD RE RE_LIO SAEB SLP_LCTRL TK VDDHD VDDI VSSI WE WE_LIO 
+ WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] 
+ WLPY_UP[3] WLP_SAE WLP_SAE_TK YL[0] YL[1] YL_LIO[0] YL_LIO[1]
*.PININFO DSLP_BUF:I SLP_LCTRL:I BLEQ_DN:O BLEQ_UP:O DEC_Y_DN[0]:O 
*.PININFO DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O DEC_Y_DN[4]:O 
*.PININFO DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O DEC_Y_UP[0]:O 
*.PININFO DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O DEC_Y_UP[4]:O 
*.PININFO DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O LIOPD:O RE_LIO:O SAEB:O 
*.PININFO WE_LIO:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B RE:B TK:B VDDHD:B VDDI:B VSSI:B WE:B WLP_SAE:B 
*.PININFO WLP_SAE_TK:B YL[0]:B YL[1]:B
XLCTRL BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ DSLP_BUF LIOPD RE RE_LIO SAEB SLP_LCTRL TK VDDHD VDDI VSSI WE WE_LIO 
+ WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] 
+ WLPY_UP[3] WLP_SAE WLP_SAE_TK YL[0] YL[1] YL_LIO[0] YL_LIO[1] S1BSVTSWSO8000Y24_LCTRL_S_M8_SD
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    XDRV_LA512_NOR_SHA
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD SLP_LCTRL TK VDDHD VDDI VSSI WE 
+ WLOUT[0] WLOUT[1] WLPY WLPYB WLP_SAE WLP_SAE_TK YL[0] YL[1]
*.PININFO DSLP_BUF:I SLP_LCTRL:I WLPY:I WLPYB:I WLP_SAE:I WLOUT[0]:O 
*.PININFO WLOUT[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B RE:B SH_NPD:B TK:B VDDHD:B VDDI:B VSSI:B WE:B 
*.PININFO WLP_SAE_TK:B YL[0]:B YL[1]:B
MM26 MWL2A MWL1A VDDI VDDI pch_mac L=35.0N W=0.5U M=2
MM23_MIXV_SLH WLOUT[1] MWL2A VDDHD VDDI pch_mac L=35.0N W=0.875U M=6
MM20_MIXV_SLH WLOUT[0] MWL2 VDDHD VDDI pch_mac L=35.0N W=0.875U M=6
MM28 MWL2A WLPY VDDI VDDI pch_mac L=35.0N W=0.64U M=2
MM18 MWL2 MWL1 VDDI VDDI pch_mac L=35.0N W=0.5U M=2
MP4 VDDHD SLP_LCTRL VDDI VDDI pch_mac L=35.0N W=0.75U M=4
MM27 MWL2 WLPY VDDI VDDI pch_mac L=35.0N W=0.64U M=2
MP6 MWL1 DEC_X0[0] SH_NPD VDDI pch_mac L=35.0N W=400N M=1
MM12 MWL1A DEC_X0[1] SH_NPD VDDI pch_mac L=35.0N W=400N M=1
MM24_MIXV_SLH WLOUT[1] MWL2A VSSI VSSI nch_mac L=35.0N W=0.65U M=4
MM15 MWL1A DEC_X0[1] VSSI VSSI nch_mac L=35.0N W=120N M=1
MM19_MIXV_SLH WLOUT[0] MWL2 VSSI VSSI nch_mac L=35.0N W=0.65U M=4
MM25 MWL2A MWL1A WLPYB VSSI nch_mac L=35.0N W=0.9U M=2
MP9 MWL1 DEC_X0[0] VSSI VSSI nch_mac L=35.0N W=120N M=1
MM6 MWL1 DEC_X1[0] VSSI VSSI nch_mac L=35.0N W=120N M=1
MM17 MWL2 MWL1 WLPYB VSSI nch_mac L=35.0N W=0.9U M=2
MM14 MWL1A DEC_X1[0] VSSI VSSI nch_mac L=35.0N W=120N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    XDRV_LA512_SHA_PMOS
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS DEC_X1 SH_NPD VDDI
*.PININFO DEC_X1:B SH_NPD:B VDDI:B
MM0 SH_NPD DEC_X1 VDDI VDDI pch_mac L=35.0N W=0.8U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    IO_M16B_WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_IO_M16B_WOBIST AWT BWEB BWEBM CKD D DM GBL GBLB GW GWB PDIO Q SLP_Q 
+ VDDF VDDFHD VDDHD VDDI VSSI WLP_SAEB
*.PININFO AWT:I BWEB:I BWEBM:I CKD:I D:I DM:I SLP_Q:I WLP_SAEB:I GW:O GWB:O 
*.PININFO Q:O GBL:B GBLB:B PDIO:B VDDF:B VDDFHD:B VDDHD:B VDDI:B VSSI:B
XIO AWT BWEB BWEBM CKD D DM GBL GBLB GW GWB Q SLP_Q VDDF VDDFHD VDDHD VDDI 
+ VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_WOBIST
MP1 VDDHD PDIO VDDI VDDI pch_mac L=35.0N W=1U M=20
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    WOBIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_WOBIST A AX VDDHD VDDI VSSI
*.PININFO A:I AX:O VDDHD:B VDDI:B VSSI:B
MM22 AX A VSSI VSSI nch_mac L=30N W=570N M=1
MM31 AX A VDDHD VDDI pch_mac L=30N W=730N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    WOBIST_WOLS_IO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_WOBIST_WOLS_IO BWEB BWEBX D DX VDDHD VDDI VSSI
*.PININFO BWEB:I D:I BWEBX:O DX:O VDDHD:B VDDI:B VSSI:B
XBIST_IO_BWEB BWEB BWEBX VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_IO_D D DX VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    REPEATER
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_REPEATER DEC0_IN[0] DEC0_IN[1] DEC0_IN[2] DEC0_IN[3] DEC0_IN[4] 
+ DEC0_IN[5] DEC0_IN[6] DEC0_IN[7] DEC0_OUT[0] DEC0_OUT[1] DEC0_OUT[2] 
+ DEC0_OUT[3] DEC0_OUT[4] DEC0_OUT[5] DEC0_OUT[6] DEC0_OUT[7] DEC1_IN[0] 
+ DEC1_IN[1] DEC1_IN[2] DEC1_IN[3] DEC1_IN[4] DEC1_IN[5] DEC1_IN[6] DEC1_IN[7] 
+ DEC1_OUT[0] DEC1_OUT[1] DEC1_OUT[2] DEC1_OUT[3] DEC1_OUT[4] DEC1_OUT[5] 
+ DEC1_OUT[6] DEC1_OUT[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DSLP_BUF RE SLP_LCTRL_IN SLP_LCTRL_OUT TK VDDHD VDDI VSSI WE WLP_SAE 
+ WLP_SAE_TK YL[0] YL[1]
*.PININFO DEC0_IN[0]:I DEC0_IN[1]:I DEC0_IN[2]:I DEC0_IN[3]:I DEC0_IN[4]:I 
*.PININFO DEC0_IN[5]:I DEC0_IN[6]:I DEC0_IN[7]:I DEC1_IN[0]:I DEC1_IN[1]:I 
*.PININFO DEC1_IN[2]:I DEC1_IN[3]:I DEC1_IN[4]:I DEC1_IN[5]:I DEC1_IN[6]:I 
*.PININFO DEC1_IN[7]:I DSLP_BUF:I SLP_LCTRL_IN:I DEC0_OUT[0]:O DEC0_OUT[1]:O 
*.PININFO DEC0_OUT[2]:O DEC0_OUT[3]:O DEC0_OUT[4]:O DEC0_OUT[5]:O 
*.PININFO DEC0_OUT[6]:O DEC0_OUT[7]:O DEC1_OUT[0]:O DEC1_OUT[1]:O 
*.PININFO DEC1_OUT[2]:O DEC1_OUT[3]:O DEC1_OUT[4]:O DEC1_OUT[5]:O 
*.PININFO DEC1_OUT[6]:O DEC1_OUT[7]:O SLP_LCTRL_OUT:O DEC_X2[0]:B DEC_X2[1]:B 
*.PININFO DEC_X2[2]:B DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B 
*.PININFO DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B 
*.PININFO DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B 
*.PININFO DEC_Y[6]:B DEC_Y[7]:B RE:B TK:B VDDHD:B VDDI:B VSSI:B WE:B WLP_SAE:B 
*.PININFO WLP_SAE_TK:B YL[0]:B YL[1]:B
XI82 NET58 VSSI VSSI VDDI VDDI SLP_LCTRL_OUT S1BSVTSWSO8000Y24_INV_BULK FN=8 WN=0.4U LN=0.03U 
+ MULTI=1 FP=8 WP=0.8U LP=0.03U
XI58[0] DEC0_IN[0] VSSI VSSI VDDI VDDI DEC0_OUT[0] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI58[1] DEC0_IN[1] VSSI VSSI VDDI VDDI DEC0_OUT[1] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI58[2] DEC0_IN[2] VSSI VSSI VDDI VDDI DEC0_OUT[2] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI58[3] DEC0_IN[3] VSSI VSSI VDDI VDDI DEC0_OUT[3] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI58[4] DEC0_IN[4] VSSI VSSI VDDI VDDI DEC0_OUT[4] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI58[5] DEC0_IN[5] VSSI VSSI VDDI VDDI DEC0_OUT[5] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI58[6] DEC0_IN[6] VSSI VSSI VDDI VDDI DEC0_OUT[6] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI58[7] DEC0_IN[7] VSSI VSSI VDDI VDDI DEC0_OUT[7] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI83 SLP_LCTRL_IN VSSI VSSI VDDI VDDI NET58 S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.4U LN=0.03U 
+ MULTI=1 FP=2 WP=0.8U LP=0.03U
XI79[0] DEC1_IN[0] VSSI VSSI VDDI VDDI DEC1_OUT[0] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI79[1] DEC1_IN[1] VSSI VSSI VDDI VDDI DEC1_OUT[1] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI79[2] DEC1_IN[2] VSSI VSSI VDDI VDDI DEC1_OUT[2] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI79[3] DEC1_IN[3] VSSI VSSI VDDI VDDI DEC1_OUT[3] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI79[4] DEC1_IN[4] VSSI VSSI VDDI VDDI DEC1_OUT[4] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI79[5] DEC1_IN[5] VSSI VSSI VDDI VDDI DEC1_OUT[5] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI79[6] DEC1_IN[6] VSSI VSSI VDDI VDDI DEC1_OUT[6] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
XI79[7] DEC1_IN[7] VSSI VSSI VDDI VDDI DEC1_OUT[7] S1BSVTSWSO8000Y24_INV_BULK FN=10 WN=0.6U 
+ LN=0.03U MULTI=1 FP=10 WP=0.6U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    YPASS_M8_16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_YPASS_M8_16 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] 
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLEQ BLEQB DL DLB READ 
+ VDDAI VDDI VSSI WC WRITE WT Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
*.PININFO BLEQ:I READ:I WRITE:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I 
*.PININFO Y[6]:I Y[7]:I BLEQB:O BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B 
*.PININFO BL[5]:B BL[6]:B BL[7]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B DL:B DLB:B VDDAI:B VDDI:B VSSI:B WC:B WT:B
XINV0 BLEQ VSSI VSSI VDDAI VDDI BLEQB S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.3U LN=0.03U MULTI=1 
+ FP=2 WP=0.95U LP=0.03U
XI246[0] YB_WRITE[0] VSSI VSSI VDDAI VDDI Y_WRITE[0] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U 
+ LN=0.03U MULTI=1 FP=1 WP=0.195U LP=0.03U
XI246[1] YB_WRITE[1] VSSI VSSI VDDAI VDDI Y_WRITE[1] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U 
+ LN=0.03U MULTI=1 FP=1 WP=0.195U LP=0.03U
XI246[2] YB_WRITE[2] VSSI VSSI VDDAI VDDI Y_WRITE[2] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U 
+ LN=0.03U MULTI=1 FP=1 WP=0.195U LP=0.03U
XI246[3] YB_WRITE[3] VSSI VSSI VDDAI VDDI Y_WRITE[3] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U 
+ LN=0.03U MULTI=1 FP=1 WP=0.195U LP=0.03U
XI246[4] YB_WRITE[4] VSSI VSSI VDDAI VDDI Y_WRITE[4] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U 
+ LN=0.03U MULTI=1 FP=1 WP=0.195U LP=0.03U
XI246[5] YB_WRITE[5] VSSI VSSI VDDAI VDDI Y_WRITE[5] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U 
+ LN=0.03U MULTI=1 FP=1 WP=0.195U LP=0.03U
XI246[6] YB_WRITE[6] VSSI VSSI VDDAI VDDI Y_WRITE[6] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U 
+ LN=0.03U MULTI=1 FP=1 WP=0.195U LP=0.03U
XI246[7] YB_WRITE[7] VSSI VSSI VDDAI VDDI Y_WRITE[7] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U 
+ LN=0.03U MULTI=1 FP=1 WP=0.195U LP=0.03U
XI244[0] Y[0] NET0116[0] VSSI VDDAI VDDI YB_READ[0] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U 
+ LN=0.03U MULTI=1 FP=1 WP=0.12U LP=0.03U
XI244[1] Y[1] NET0116[1] VSSI VDDAI VDDI YB_READ[1] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U 
+ LN=0.03U MULTI=1 FP=1 WP=0.12U LP=0.03U
XI244[2] Y[2] NET0116[2] VSSI VDDAI VDDI YB_READ[2] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U 
+ LN=0.03U MULTI=1 FP=1 WP=0.12U LP=0.03U
XI244[3] Y[3] NET0116[3] VSSI VDDAI VDDI YB_READ[3] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U 
+ LN=0.03U MULTI=1 FP=1 WP=0.12U LP=0.03U
XI244[4] Y[4] NET0116[4] VSSI VDDAI VDDI YB_READ[4] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U 
+ LN=0.03U MULTI=1 FP=1 WP=0.12U LP=0.03U
XI244[5] Y[5] NET0116[5] VSSI VDDAI VDDI YB_READ[5] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U 
+ LN=0.03U MULTI=1 FP=1 WP=0.12U LP=0.03U
XI244[6] Y[6] NET0116[6] VSSI VDDAI VDDI YB_READ[6] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U 
+ LN=0.03U MULTI=1 FP=1 WP=0.12U LP=0.03U
XI244[7] Y[7] NET0116[7] VSSI VDDAI VDDI YB_READ[7] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U 
+ LN=0.03U MULTI=1 FP=1 WP=0.12U LP=0.03U
XI245[0] Y[0] NET0112[0] VSSI VDDAI VDDI YB_WRITE[0] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.20U 
+ LN=0.03U MULTI=1 FP=1 WP=0.15U LP=0.03U
XI245[1] Y[1] NET0112[1] VSSI VDDAI VDDI YB_WRITE[1] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.20U 
+ LN=0.03U MULTI=1 FP=1 WP=0.15U LP=0.03U
XI245[2] Y[2] NET0112[2] VSSI VDDAI VDDI YB_WRITE[2] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.20U 
+ LN=0.03U MULTI=1 FP=1 WP=0.15U LP=0.03U
XI245[3] Y[3] NET0112[3] VSSI VDDAI VDDI YB_WRITE[3] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.20U 
+ LN=0.03U MULTI=1 FP=1 WP=0.15U LP=0.03U
XI245[4] Y[4] NET0112[4] VSSI VDDAI VDDI YB_WRITE[4] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.20U 
+ LN=0.03U MULTI=1 FP=1 WP=0.15U LP=0.03U
XI245[5] Y[5] NET0112[5] VSSI VDDAI VDDI YB_WRITE[5] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.20U 
+ LN=0.03U MULTI=1 FP=1 WP=0.15U LP=0.03U
XI245[6] Y[6] NET0112[6] VSSI VDDAI VDDI YB_WRITE[6] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.20U 
+ LN=0.03U MULTI=1 FP=1 WP=0.15U LP=0.03U
XI245[7] Y[7] NET0112[7] VSSI VDDAI VDDI YB_WRITE[7] S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.20U 
+ LN=0.03U MULTI=1 FP=1 WP=0.15U LP=0.03U
MP17[0] YB_READ[0] READ VDDAI VDDI pch_mac L=30N W=120N M=1
MP17[1] YB_READ[1] READ VDDAI VDDI pch_mac L=30N W=120N M=1
MP17[2] YB_READ[2] READ VDDAI VDDI pch_mac L=30N W=120N M=1
MP17[3] YB_READ[3] READ VDDAI VDDI pch_mac L=30N W=120N M=1
MP17[4] YB_READ[4] READ VDDAI VDDI pch_mac L=30N W=120N M=1
MP17[5] YB_READ[5] READ VDDAI VDDI pch_mac L=30N W=120N M=1
MP17[6] YB_READ[6] READ VDDAI VDDI pch_mac L=30N W=120N M=1
MP17[7] YB_READ[7] READ VDDAI VDDI pch_mac L=30N W=120N M=1
MP10_MIXV_SLS[0] DLB YB_READ[0] BLB[0] VDDI pch_mac L=30N W=370N M=1
MP10_MIXV_SLS[1] DLB YB_READ[1] BLB[1] VDDI pch_mac L=30N W=370N M=1
MP10_MIXV_SLS[2] DLB YB_READ[2] BLB[2] VDDI pch_mac L=30N W=370N M=1
MP10_MIXV_SLS[3] DLB YB_READ[3] BLB[3] VDDI pch_mac L=30N W=370N M=1
MP10_MIXV_SLS[4] DLB YB_READ[4] BLB[4] VDDI pch_mac L=30N W=370N M=1
MP10_MIXV_SLS[5] DLB YB_READ[5] BLB[5] VDDI pch_mac L=30N W=370N M=1
MP10_MIXV_SLS[6] DLB YB_READ[6] BLB[6] VDDI pch_mac L=30N W=370N M=1
MP10_MIXV_SLS[7] DLB YB_READ[7] BLB[7] VDDI pch_mac L=30N W=370N M=1
MP3 DLB BLEQB VDDAI VDDI pch_mac L=30N W=120N M=1
MP0_MIXV_SLS[0] DL YB_READ[0] BL[0] VDDI pch_mac L=30N W=370N M=1
MP0_MIXV_SLS[1] DL YB_READ[1] BL[1] VDDI pch_mac L=30N W=370N M=1
MP0_MIXV_SLS[2] DL YB_READ[2] BL[2] VDDI pch_mac L=30N W=370N M=1
MP0_MIXV_SLS[3] DL YB_READ[3] BL[3] VDDI pch_mac L=30N W=370N M=1
MP0_MIXV_SLS[4] DL YB_READ[4] BL[4] VDDI pch_mac L=30N W=370N M=1
MP0_MIXV_SLS[5] DL YB_READ[5] BL[5] VDDI pch_mac L=30N W=370N M=1
MP0_MIXV_SLS[6] DL YB_READ[6] BL[6] VDDI pch_mac L=30N W=370N M=1
MP0_MIXV_SLS[7] DL YB_READ[7] BL[7] VDDI pch_mac L=30N W=370N M=1
MP22 VDDAI BLEQB DL VDDI pch_mac L=30N W=120N M=1
MP29[0] YB_WRITE[0] WRITE VDDAI VDDI pch_mac L=30N W=150N M=1
MP29[1] YB_WRITE[1] WRITE VDDAI VDDI pch_mac L=30N W=150N M=1
MP29[2] YB_WRITE[2] WRITE VDDAI VDDI pch_mac L=30N W=150N M=1
MP29[3] YB_WRITE[3] WRITE VDDAI VDDI pch_mac L=30N W=150N M=1
MP29[4] YB_WRITE[4] WRITE VDDAI VDDI pch_mac L=30N W=150N M=1
MP29[5] YB_WRITE[5] WRITE VDDAI VDDI pch_mac L=30N W=150N M=1
MP29[6] YB_WRITE[6] WRITE VDDAI VDDI pch_mac L=30N W=150N M=1
MP29[7] YB_WRITE[7] WRITE VDDAI VDDI pch_mac L=30N W=150N M=1
MM3_MIXV_SLH[0] BL[0] BLB[0] VDDAI VDDI pch_mac L=30N W=120N M=1
MM3_MIXV_SLH[1] BL[1] BLB[1] VDDAI VDDI pch_mac L=30N W=120N M=1
MM3_MIXV_SLH[2] BL[2] BLB[2] VDDAI VDDI pch_mac L=30N W=120N M=1
MM3_MIXV_SLH[3] BL[3] BLB[3] VDDAI VDDI pch_mac L=30N W=120N M=1
MM3_MIXV_SLH[4] BL[4] BLB[4] VDDAI VDDI pch_mac L=30N W=120N M=1
MM3_MIXV_SLH[5] BL[5] BLB[5] VDDAI VDDI pch_mac L=30N W=120N M=1
MM3_MIXV_SLH[6] BL[6] BLB[6] VDDAI VDDI pch_mac L=30N W=120N M=1
MM3_MIXV_SLH[7] BL[7] BLB[7] VDDAI VDDI pch_mac L=30N W=120N M=1
MM2_MIXV_SLH[0] BLB[0] BL[0] VDDAI VDDI pch_mac L=30N W=120N M=1
MM2_MIXV_SLH[1] BLB[1] BL[1] VDDAI VDDI pch_mac L=30N W=120N M=1
MM2_MIXV_SLH[2] BLB[2] BL[2] VDDAI VDDI pch_mac L=30N W=120N M=1
MM2_MIXV_SLH[3] BLB[3] BL[3] VDDAI VDDI pch_mac L=30N W=120N M=1
MM2_MIXV_SLH[4] BLB[4] BL[4] VDDAI VDDI pch_mac L=30N W=120N M=1
MM2_MIXV_SLH[5] BLB[5] BL[5] VDDAI VDDI pch_mac L=30N W=120N M=1
MM2_MIXV_SLH[6] BLB[6] BL[6] VDDAI VDDI pch_mac L=30N W=120N M=1
MM2_MIXV_SLH[7] BLB[7] BL[7] VDDAI VDDI pch_mac L=30N W=120N M=1
MN31_MIXV_SLS[0] BL[0] Y_WRITE[0] WT VSSI nch_mac L=30N W=850N M=1
MN31_MIXV_SLS[1] BL[1] Y_WRITE[1] WT VSSI nch_mac L=30N W=850N M=1
MN31_MIXV_SLS[2] BL[2] Y_WRITE[2] WT VSSI nch_mac L=30N W=850N M=1
MN31_MIXV_SLS[3] BL[3] Y_WRITE[3] WT VSSI nch_mac L=30N W=850N M=1
MN31_MIXV_SLS[4] BL[4] Y_WRITE[4] WT VSSI nch_mac L=30N W=850N M=1
MN31_MIXV_SLS[5] BL[5] Y_WRITE[5] WT VSSI nch_mac L=30N W=850N M=1
MN31_MIXV_SLS[6] BL[6] Y_WRITE[6] WT VSSI nch_mac L=30N W=850N M=1
MN31_MIXV_SLS[7] BL[7] Y_WRITE[7] WT VSSI nch_mac L=30N W=850N M=1
MN18_MIXV_SLS[0] BLB[0] Y_WRITE[0] WC VSSI nch_mac L=30N W=850N M=1
MN18_MIXV_SLS[1] BLB[1] Y_WRITE[1] WC VSSI nch_mac L=30N W=850N M=1
MN18_MIXV_SLS[2] BLB[2] Y_WRITE[2] WC VSSI nch_mac L=30N W=850N M=1
MN18_MIXV_SLS[3] BLB[3] Y_WRITE[3] WC VSSI nch_mac L=30N W=850N M=1
MN18_MIXV_SLS[4] BLB[4] Y_WRITE[4] WC VSSI nch_mac L=30N W=850N M=1
MN18_MIXV_SLS[5] BLB[5] Y_WRITE[5] WC VSSI nch_mac L=30N W=850N M=1
MN18_MIXV_SLS[6] BLB[6] Y_WRITE[6] WC VSSI nch_mac L=30N W=850N M=1
MN18_MIXV_SLS[7] BLB[7] Y_WRITE[7] WC VSSI nch_mac L=30N W=850N M=1
MN13[0] NET0116[0] READ VSSI VSSI nch_mac L=30N W=310N M=1
MN13[1] NET0116[1] READ VSSI VSSI nch_mac L=30N W=310N M=1
MN13[2] NET0116[2] READ VSSI VSSI nch_mac L=30N W=310N M=1
MN13[3] NET0116[3] READ VSSI VSSI nch_mac L=30N W=310N M=1
MN13[4] NET0116[4] READ VSSI VSSI nch_mac L=30N W=310N M=1
MN13[5] NET0116[5] READ VSSI VSSI nch_mac L=30N W=310N M=1
MN13[6] NET0116[6] READ VSSI VSSI nch_mac L=30N W=310N M=1
MN13[7] NET0116[7] READ VSSI VSSI nch_mac L=30N W=310N M=1
MN1[0] NET0112[0] WRITE VSSI VSSI nch_mac L=30N W=310N M=1
MN1[1] NET0112[1] WRITE VSSI VSSI nch_mac L=30N W=310N M=1
MN1[2] NET0112[2] WRITE VSSI VSSI nch_mac L=30N W=310N M=1
MN1[3] NET0112[3] WRITE VSSI VSSI nch_mac L=30N W=310N M=1
MN1[4] NET0112[4] WRITE VSSI VSSI nch_mac L=30N W=310N M=1
MN1[5] NET0112[5] WRITE VSSI VSSI nch_mac L=30N W=310N M=1
MN1[6] NET0112[6] WRITE VSSI VSSI nch_mac L=30N W=310N M=1
MN1[7] NET0112[7] WRITE VSSI VSSI nch_mac L=30N W=310N M=1
XPRECHARGE[0] BL[0] BLB[0] BLEQB VDDAI VDDI S1BSVTSWSO8000Y24_PRECHARGE
XPRECHARGE[1] BL[1] BLB[1] BLEQB VDDAI VDDI S1BSVTSWSO8000Y24_PRECHARGE
XPRECHARGE[2] BL[2] BLB[2] BLEQB VDDAI VDDI S1BSVTSWSO8000Y24_PRECHARGE
XPRECHARGE[3] BL[3] BLB[3] BLEQB VDDAI VDDI S1BSVTSWSO8000Y24_PRECHARGE
XPRECHARGE[4] BL[4] BLB[4] BLEQB VDDAI VDDI S1BSVTSWSO8000Y24_PRECHARGE
XPRECHARGE[5] BL[5] BLB[5] BLEQB VDDAI VDDI S1BSVTSWSO8000Y24_PRECHARGE
XPRECHARGE[6] BL[6] BLB[6] BLEQB VDDAI VDDI S1BSVTSWSO8000Y24_PRECHARGE
XPRECHARGE[7] BL[7] BLB[7] BLEQB VDDAI VDDI S1BSVTSWSO8000Y24_PRECHARGE
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    SA_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_SA_M16 DLB_DN_0 DLB_DN_1 DLB_UP_0 DLB_UP_1 DL_DN_0 DL_DN_1 DL_UP_0 
+ DL_UP_1 GBL GBLB PGB_DN_0 PGB_DN_1 PGB_UP_0 PGB_UP_1 PREB SAE VDDAI VDDI VSSI
*.PININFO PGB_DN_0:I PGB_DN_1:I PGB_UP_0:I PGB_UP_1:I PREB:I SAE:I DLB_DN_0:B 
*.PININFO DLB_DN_1:B DLB_UP_0:B DLB_UP_1:B DL_DN_0:B DL_DN_1:B DL_UP_0:B 
*.PININFO DL_UP_1:B GBL:B GBLB:B VDDAI:B VDDI:B VSSI:B
MN0 DL_IN DLB_IN NS VSSI nch_mac L=90N W=0.5U M=4
MN2 NS SAE VSSI VSSI nch_mac L=30N W=0.5U M=4
MN1 DLB_IN DL_IN NS VSSI nch_mac L=90N W=0.5U M=4
MN11 GBL SO VSSI VSSI nch_mac L=35.0N W=0.95U M=3
MN12 GBLB SOB VSSI VSSI nch_mac L=35.0N W=0.95U M=3
MP2 DL_IN DLB_IN VDDAI VDDI pch_mac L=30N W=500N M=1
MP10 DL_IN PREB VDDAI VDDI pch_mac L=30N W=500N M=1
MP6 DL_UP_0 PGB_UP_0 DL_IN VDDI pch_mac L=30N W=500N M=1
MP0 DLB_UP_1 PGB_UP_1 DLB_IN VDDI pch_mac L=30N W=500N M=1
MP7 DLB_UP_0 PGB_UP_0 DLB_IN VDDI pch_mac L=30N W=500N M=1
MP13 DL_DN_1 PGB_DN_1 DL_IN VDDI pch_mac L=30N W=500N M=1
MP3 DLB_IN DL_IN VDDAI VDDI pch_mac L=30N W=500N M=1
MP14 DLB_DN_1 PGB_DN_1 DLB_IN VDDI pch_mac L=30N W=500N M=1
MP8 DL_IN PREB DLB_IN VDDI pch_mac L=30N W=0.5U M=2
MP11 DLB_IN PREB VDDAI VDDI pch_mac L=30N W=500N M=1
MP4 DL_DN_0 PGB_DN_0 DL_IN VDDI pch_mac L=30N W=500N M=1
MP1 DL_UP_1 PGB_UP_1 DL_IN VDDI pch_mac L=30N W=500N M=1
MP5 DLB_DN_0 PGB_DN_0 DLB_IN VDDI pch_mac L=30N W=500N M=1
XINV0 DL_IN VSSI VSSI VDDAI VDDI SO S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U LN=0.03U MULTI=1 
+ FP=3 WP=0.22U LP=0.03U
XINV1 DLB_IN VSSI VSSI VDDAI VDDI SOB S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.2U LN=0.03U MULTI=1 
+ FP=3 WP=0.22U LP=0.03U
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    IO_RWBLK_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_IO_RWBLK_M16 BLEQB_DN_0 BLEQB_DN_1 BLEQB_UP_0 BLEQB_UP_1 BLEQ_DN 
+ BLEQ_UP DLB_DN_0 DLB_DN_1 DLB_UP_0 DLB_UP_1 DL_DN_0 DL_DN_1 DL_UP_0 DL_UP_1 
+ GBL GBLB GW GWB RE READ SAEB VDDAI VDDI VSSI WC[0] WC[1] WE WRITE WT[0] 
+ WT[1] YL[0] YL[1]
*.PININFO BLEQB_DN_0:I BLEQB_DN_1:I BLEQB_UP_0:I BLEQB_UP_1:I BLEQ_DN:I 
*.PININFO BLEQ_UP:I GW:I GWB:I RE:I SAEB:I WE:I YL[0]:I YL[1]:I READ:O WC[0]:O 
*.PININFO WC[1]:O WRITE:O WT[0]:O WT[1]:O DLB_DN_0:B DLB_DN_1:B DLB_UP_0:B 
*.PININFO DLB_UP_1:B DL_DN_0:B DL_DN_1:B DL_UP_0:B DL_UP_1:B GBL:B GBLB:B 
*.PININFO VDDAI:B VDDI:B VSSI:B
XI100 BLEQ_UP VSSI VSSI VDDAI VDDI NET0227 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XI99 BLEQ_DN VSSI VSSI VDDAI VDDI NET0228 S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XI1 WE VSSI VSSI VDDAI VDDI WE1B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.24U LP=0.03U
XI97 NET0228 VSSI VSSI VDDAI VDDI BLEQ2_DN S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XI96 NET0227 VSSI VSSI VDDAI VDDI BLEQ2_UP S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U 
+ MULTI=1 FP=1 WP=0.12U LP=0.03U
XINV4 WE1B VSSI VSSI VDDAI VDDI WRITE S1BSVTSWSO8000Y24_INV_BULK FN=5 WN=0.2U LN=0.03U MULTI=1 
+ FP=5 WP=0.5U LP=0.03U
XINV5 RE1B VSSI VSSI VDDAI VDDI READ S1BSVTSWSO8000Y24_INV_BULK FN=5 WN=0.2U LN=0.03U MULTI=1 
+ FP=5 WP=0.5U LP=0.03U
XI248 SAEC VSSI VSSI VDDAI VDDI SAE S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.3U LP=0.03U
XI2 RE VSSI VSSI VDDAI VDDI RE1B S1BSVTSWSO8000Y24_INV_BULK FN=1 WN=0.12U LN=0.03U MULTI=1 
+ FP=1 WP=0.24U LP=0.03U
XI89 GWDC_YLB VSSI VSSI VDDAI VDDI LWDC[0] S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.2U LN=0.03U 
+ MULTI=1 FP=2 WP=0.3U LP=0.03U
XI90 GWDT_YLB VSSI VSSI VDDAI VDDI LWDT[0] S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.2U LN=0.03U 
+ MULTI=1 FP=2 WP=0.3U LP=0.03U
XI91 GWDT_YL VSSI VSSI VDDAI VDDI LWDT[1] S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.2U LN=0.03U 
+ MULTI=1 FP=2 WP=0.3U LP=0.03U
XI88 GWDC_YL VSSI VSSI VDDAI VDDI LWDC[1] S1BSVTSWSO8000Y24_INV_BULK FN=2 WN=0.2U LN=0.03U 
+ MULTI=1 FP=2 WP=0.3U LP=0.03U
XI76 BLEQB_UP_1 YL[1] VSSI VSSI VDDAI VDDI PGB_UP_1 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.2U 
+ LN1=0.03U FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.3U LP1=0.03U
XI78 BLEQB_DN_1 YL[1] VSSI VSSI VDDAI VDDI PGB_DN_1 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.2U 
+ LN1=0.03U FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.3U LP1=0.03U
XI77 BLEQB_DN_0 YL[0] VSSI VSSI VDDAI VDDI PGB_DN_0 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.2U 
+ LN1=0.03U FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.3U LP1=0.03U
XI75 BLEQB_UP_0 YL[0] VSSI VSSI VDDAI VDDI PGB_UP_0 S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.2U 
+ LN1=0.03U FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.3U LP1=0.03U
XI92 GW YL[0] VSSI VSSI VDDAI VDDI GWDT_YLB S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.2U 
+ LN1=0.03U FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.3U LP1=0.03U
XI94 GWB YL[0] VSSI VSSI VDDAI VDDI GWDC_YLB S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.2U 
+ LN1=0.03U FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.3U LP1=0.03U
XI93 GW YL[1] VSSI VSSI VDDAI VDDI GWDT_YL S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.2U 
+ LN1=0.03U FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.3U LP1=0.03U
XI28 GWB YL[1] VSSI VSSI VDDAI VDDI GWDC_YL S1BSVTSWSO8000Y24_NAND_BULK FN1=1 WN1=0.2U 
+ LN1=0.03U FN2=1 WN2=0.2U LN2=0.03U FP2=1 WP2=0.3U LP2=0.03U MULTI=1 FP1=1 
+ WP1=0.3U LP1=0.03U
XI222 SAEC BLEQ2_UP BLEQ2_DN VSSI VSSI VDDAI VDDI PREB S1BSVTSWSO8000Y24_NAND3_BULK FN1=1 
+ WN1=0.3U LN1=0.03U FN2=1 WN2=0.3U LN2=0.03U FN3=1 WN3=0.3U LN3=0.03U FP3=1 
+ WP3=0.2U LP3=0.03U FP2=1 WP2=0.2U LP2=0.03U MULTI=1 FP1=1 WP1=0.2U LP1=0.03U
XI235 GBLB GBL SAEB VSSI VSSI VDDAI VDDI SAEC S1BSVTSWSO8000Y24_NAND3_BULK FN1=1 WN1=0.29U 
+ LN1=0.03U FN2=1 WN2=0.29U LN2=0.03U FN3=1 WN3=0.29U LN3=0.03U FP3=1 WP3=0.2U 
+ LP3=0.03U FP2=1 WP2=0.2U LP2=0.03U MULTI=1 FP1=1 WP1=0.2U LP1=0.03U
MN0 WC[1] LWDT[1] VSSI VSSI nch_mac L=30N W=0.57U M=6
MM4 WT[0] LWDC[0] VSSI VSSI nch_mac L=30N W=0.57U M=6
MM3 WT[1] LWDC[1] VSSI VSSI nch_mac L=30N W=0.57U M=6
MM0 WC[0] LWDT[0] VSSI VSSI nch_mac L=30N W=0.57U M=6
MP27 WC[1] LWDT[1] VDDAI VDDI pch_mac L=30N W=0.56U M=2
MM2 WT[1] LWDC[1] VDDAI VDDI pch_mac L=30N W=0.56U M=2
MM1 WC[0] LWDT[0] VDDAI VDDI pch_mac L=30N W=0.56U M=2
MM5 WT[0] LWDC[0] VDDAI VDDI pch_mac L=30N W=0.56U M=2
XSA DLB_DN_0 DLB_DN_1 DLB_UP_0 DLB_UP_1 DL_DN_0 DL_DN_1 DL_UP_0 DL_UP_1 GBL 
+ GBLB PGB_DN_0 PGB_DN_1 PGB_UP_0 PGB_UP_1 PREB SAE VDDAI VDDI VSSI S1BSVTSWSO8000Y24_SA_M16
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    LIO_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_LIO_M16 BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12] 
+ BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] 
+ BLB_UP[4] BLB_UP[5] BLB_UP[6] BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10] 
+ BLB_UP[11] BLB_UP[12] BLB_UP[13] BLB_UP[14] BLB_UP[15] BLEQ_DN BLEQ_UP 
+ BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] 
+ BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14] 
+ BL_DN[15] BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] 
+ BL_UP[7] BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14] 
+ BL_UP[15] GBL GBLB GW GWB RE SAEB VDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] 
+ Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] 
+ Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
*.PININFO BLEQ_DN:I BLEQ_UP:I GW:I GWB:I RE:I SAEB:I WE:I YL_LIO[0]:I 
*.PININFO YL_LIO[1]:I Y_DN[0]:I Y_DN[1]:I Y_DN[2]:I Y_DN[3]:I Y_DN[4]:I 
*.PININFO Y_DN[5]:I Y_DN[6]:I Y_DN[7]:I Y_UP[0]:I Y_UP[1]:I Y_UP[2]:I 
*.PININFO Y_UP[3]:I Y_UP[4]:I Y_UP[5]:I Y_UP[6]:I Y_UP[7]:I BLB_DN[0]:B 
*.PININFO BLB_DN[1]:B BLB_DN[2]:B BLB_DN[3]:B BLB_DN[4]:B BLB_DN[5]:B 
*.PININFO BLB_DN[6]:B BLB_DN[7]:B BLB_DN[8]:B BLB_DN[9]:B BLB_DN[10]:B 
*.PININFO BLB_DN[11]:B BLB_DN[12]:B BLB_DN[13]:B BLB_DN[14]:B BLB_DN[15]:B 
*.PININFO BLB_UP[0]:B BLB_UP[1]:B BLB_UP[2]:B BLB_UP[3]:B BLB_UP[4]:B 
*.PININFO BLB_UP[5]:B BLB_UP[6]:B BLB_UP[7]:B BLB_UP[8]:B BLB_UP[9]:B 
*.PININFO BLB_UP[10]:B BLB_UP[11]:B BLB_UP[12]:B BLB_UP[13]:B BLB_UP[14]:B 
*.PININFO BLB_UP[15]:B BL_DN[0]:B BL_DN[1]:B BL_DN[2]:B BL_DN[3]:B BL_DN[4]:B 
*.PININFO BL_DN[5]:B BL_DN[6]:B BL_DN[7]:B BL_DN[8]:B BL_DN[9]:B BL_DN[10]:B 
*.PININFO BL_DN[11]:B BL_DN[12]:B BL_DN[13]:B BL_DN[14]:B BL_DN[15]:B 
*.PININFO BL_UP[0]:B BL_UP[1]:B BL_UP[2]:B BL_UP[3]:B BL_UP[4]:B BL_UP[5]:B 
*.PININFO BL_UP[6]:B BL_UP[7]:B BL_UP[8]:B BL_UP[9]:B BL_UP[10]:B BL_UP[11]:B 
*.PININFO BL_UP[12]:B BL_UP[13]:B BL_UP[14]:B BL_UP[15]:B GBL:B GBLB:B VDDAI:B 
*.PININFO VDDI:B VSSI:B
XYPASS_UP_1 BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] 
+ BL_UP[14] BL_UP[15] BLB_UP[8] BLB_UP[9] BLB_UP[10] BLB_UP[11] BLB_UP[12] 
+ BLB_UP[13] BLB_UP[14] BLB_UP[15] BLEQ_UP BLEQB_UP_1 DL_UP_1 DLB_UP_1 READ 
+ VDDAI VDDI VSSI WC[1] WRITE WT[1] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] 
+ Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_YPASS_M8_16
XYPASS_UP_0 BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] 
+ BL_UP[7] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] BLB_UP[4] BLB_UP[5] 
+ BLB_UP[6] BLB_UP[7] BLEQ_UP BLEQB_UP_0 DL_UP_0 DLB_UP_0 READ VDDAI VDDI VSSI 
+ WC[0] WRITE WT[0] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] 
+ Y_UP[7] S1BSVTSWSO8000Y24_YPASS_M8_16
XYPASS_DN_0 BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] 
+ BL_DN[7] BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLEQ_DN BLEQB_DN_0 DL_DN_0 DLB_DN_0 READ VDDAI VDDI VSSI 
+ WC[0] WRITE WT[0] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] 
+ Y_DN[7] S1BSVTSWSO8000Y24_YPASS_M8_16
XYPASS_DN_1 BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] 
+ BL_DN[14] BL_DN[15] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12] 
+ BLB_DN[13] BLB_DN[14] BLB_DN[15] BLEQ_DN BLEQB_DN_1 DL_DN_1 DLB_DN_1 READ 
+ VDDAI VDDI VSSI WC[1] WRITE WT[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] 
+ Y_DN[5] Y_DN[6] Y_DN[7] S1BSVTSWSO8000Y24_YPASS_M8_16
XIO_RWBLK BLEQB_DN_0 BLEQB_DN_1 BLEQB_UP_0 BLEQB_UP_1 BLEQ_DN BLEQ_UP DLB_DN_0 
+ DLB_DN_1 DLB_UP_0 DLB_UP_1 DL_DN_0 DL_DN_1 DL_UP_0 DL_UP_1 GBL GBLB GW GWB 
+ RE READ SAEB VDDAI VDDI VSSI WC[0] WC[1] WE WRITE WT[0] WT[1] YL_LIO[0] 
+ YL_LIO[1] S1BSVTSWSO8000Y24_IO_RWBLK_M16
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    LIO_M16_SD
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_LIO_M16_SD BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12] 
+ BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] 
+ BLB_UP[4] BLB_UP[5] BLB_UP[6] BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10] 
+ BLB_UP[11] BLB_UP[12] BLB_UP[13] BLB_UP[14] BLB_UP[15] BLEQ_DN BLEQ_UP 
+ BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] 
+ BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14] 
+ BL_DN[15] BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] 
+ BL_UP[7] BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14] 
+ BL_UP[15] GBL GBLB GW GWB LIOPD PDI PDO PDO_BACK RE SAEB VDDAI VDDI VSSI WE 
+ YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] 
+ Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
*.PININFO BLEQ_DN:I BLEQ_UP:I GW:I GWB:I LIOPD:I PDI:I PDO_BACK:I RE:I SAEB:I 
*.PININFO WE:I YL_LIO[0]:I YL_LIO[1]:I Y_DN[0]:I Y_DN[1]:I Y_DN[2]:I Y_DN[3]:I 
*.PININFO Y_DN[4]:I Y_DN[5]:I Y_DN[6]:I Y_DN[7]:I Y_UP[0]:I Y_UP[1]:I 
*.PININFO Y_UP[2]:I Y_UP[3]:I Y_UP[4]:I Y_UP[5]:I Y_UP[6]:I Y_UP[7]:I PDO:O 
*.PININFO BLB_DN[0]:B BLB_DN[1]:B BLB_DN[2]:B BLB_DN[3]:B BLB_DN[4]:B 
*.PININFO BLB_DN[5]:B BLB_DN[6]:B BLB_DN[7]:B BLB_DN[8]:B BLB_DN[9]:B 
*.PININFO BLB_DN[10]:B BLB_DN[11]:B BLB_DN[12]:B BLB_DN[13]:B BLB_DN[14]:B 
*.PININFO BLB_DN[15]:B BLB_UP[0]:B BLB_UP[1]:B BLB_UP[2]:B BLB_UP[3]:B 
*.PININFO BLB_UP[4]:B BLB_UP[5]:B BLB_UP[6]:B BLB_UP[7]:B BLB_UP[8]:B 
*.PININFO BLB_UP[9]:B BLB_UP[10]:B BLB_UP[11]:B BLB_UP[12]:B BLB_UP[13]:B 
*.PININFO BLB_UP[14]:B BLB_UP[15]:B BL_DN[0]:B BL_DN[1]:B BL_DN[2]:B 
*.PININFO BL_DN[3]:B BL_DN[4]:B BL_DN[5]:B BL_DN[6]:B BL_DN[7]:B BL_DN[8]:B 
*.PININFO BL_DN[9]:B BL_DN[10]:B BL_DN[11]:B BL_DN[12]:B BL_DN[13]:B 
*.PININFO BL_DN[14]:B BL_DN[15]:B BL_UP[0]:B BL_UP[1]:B BL_UP[2]:B BL_UP[3]:B 
*.PININFO BL_UP[4]:B BL_UP[5]:B BL_UP[6]:B BL_UP[7]:B BL_UP[8]:B BL_UP[9]:B 
*.PININFO BL_UP[10]:B BL_UP[11]:B BL_UP[12]:B BL_UP[13]:B BL_UP[14]:B 
*.PININFO BL_UP[15]:B GBL:B GBLB:B VDDAI:B VDDI:B VSSI:B
XLIO_HEADER[0] LIOPD PDI PDO0 PDO_BACK VDDAI VDDI VSSI S1BSVTSWSO8000Y24_LIO_HEADER_N1
XLIO_HEADER[1] LIOPD PDO0 PDO1 PDO1 VDDAI VDDI VSSI S1BSVTSWSO8000Y24_LIO_HEADER_N1
XLIO_HEADER[2] LIOPD PDO1 PDO2 PDO_BACK VDDAI VDDI VSSI S1BSVTSWSO8000Y24_LIO_HEADER_N1
XLIO_HEADER[3] LIOPD PDO2 PDO3 PDO3 VDDAI VDDI VSSI S1BSVTSWSO8000Y24_LIO_HEADER_N1
XLIO_HEADER[4] LIOPD PDO3 PDO4 PDO_BACK VDDAI VDDI VSSI S1BSVTSWSO8000Y24_LIO_HEADER_N1
XLIO_HEADER[5] LIOPD PDO4 PDO5 PDO5 VDDAI VDDI VSSI S1BSVTSWSO8000Y24_LIO_HEADER_N1
XLIO_HEADER[6] LIOPD PDO5 PDO6 PDO_BACK VDDAI VDDI VSSI S1BSVTSWSO8000Y24_LIO_HEADER_N1
XLIO_HEADER[7] LIOPD PDO6 PDO PDO VDDAI VDDI VSSI S1BSVTSWSO8000Y24_LIO_HEADER_N1
XLIO BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] BLB_DN[6] 
+ BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12] BLB_DN[13] 
+ BLB_DN[14] BLB_DN[15] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] BLB_UP[4] 
+ BLB_UP[5] BLB_UP[6] BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10] BLB_UP[11] 
+ BLB_UP[12] BLB_UP[13] BLB_UP[14] BLB_UP[15] BLEQ_DN BLEQ_UP BL_DN[0] 
+ BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] BL_DN[8] 
+ BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14] BL_DN[15] 
+ BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] BL_UP[7] 
+ BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14] 
+ BL_UP[15] GBL GBLB GW GWB RE SAEB VDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] 
+ Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] 
+ Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    CLK_BUF
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_CLK_BUF IN OUT VDDHD VDDI VSSI
*.PININFO IN:I OUT:O VDDHD:B VDDI:B VSSI:B
MP3_MIXV_SLS NET66 IN VDDHD VDDI pch_mac L=30N W=300N M=1
MM2_MIXV_SLS OUT NET66 VDDHD VDDI pch_mac L=30N W=0.7U M=2
MN1_MIXV_SLS NET66 IN VSSI VSSI nch_mac L=30N W=480N M=1
MM3_MIXV_SLS OUT NET66 VSSI VSSI nch_mac L=30N W=700N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    BIST_VHILO_M8_WOWO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_BIST_VHILO_M8_WOWO VDDI VHI VLO VSSI
*.PININFO VHI:O VLO:O VDDI:B VSSI:B
MN3 VSSI Z2 Z1 VSSI nch_mac L=30N W=360N M=1
MN0 VSSI Z1 Z1 VSSI nch_mac L=30N W=360N M=1
MN1 VSSI Z2 VLO VSSI nch_mac L=30N W=0.75U M=4
MP7 Z2 Z1 VDDI VDDI pch_mac L=30N W=360N M=1
MP2 VHI Z1 VDDI VDDI pch_mac L=30N W=0.75U M=4
MP0 Z2 Z2 VDDI VDDI pch_mac L=30N W=360N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    TOP_EDGE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_TOP_EDGE VDDHD VDDI VSSI WLP_SAE WLP_SAE_TK
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
MM5 NET17 WLP_SAE VSSI VSSI nch_mac L=30N W=0.95U M=6
MM2 NET17 WLP_SAE VSSI VSSI nch_mac L=30N W=1.25U M=2
MM1 NET17 WLP_SAE VSSI VSSI nch_mac L=30N W=800N M=1
MM7 WLP_SAE_TK NET17 VSSI VSSI nch_mac L=30N W=0.65U M=6
MM12 WLP_SAE_TK NET17 VDDHD VDDI pch_mac L=30N W=0.5U M=3
MM4 WLP_SAE_TK NET17 VDDHD VDDI pch_mac L=30N W=0.9U M=3
MM11 WLP_SAE_TK NET17 VDDHD VDDI pch_mac L=30N W=0.75U M=4
MM0 NET17 WLP_SAE VDDHD VDDI pch_mac L=30N W=0.565U M=3
MM3 WLP_SAE_TK NET17 VDDHD VDDI pch_mac L=30N W=0.875U M=12
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    IO_M16B_WOBIST_SR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR AWT BWEB CKD D GBL GBLB GW GWB IOPD Q SLP_Q VDDHD 
+ VDDI VSSI WLP_SAEB
*.PININFO AWT:I BWEB:I CKD:I D:I SLP_Q:I WLP_SAEB:I GW:O GWB:O Q:O GBL:B 
*.PININFO GBLB:B IOPD:B VDDHD:B VDDI:B VSSI:B
XIO_LL AWT BWEBX NET025 CKD DX NET026 GBL GBLB GW GWB IOPD Q SLP_Q VDDI VDDHD 
+ VDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST
XIO_PAD_LL BWEB BWEBX D DX VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST_WOLS_IO
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    WOBIST_WOLS_CNT_M16_IOX2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_WOBIST_WOLS_CNT_M16_IOX2 BWEBX_L BWEBX_R BWEB_L BWEB_R CEB CEB3B CLK 
+ CLK2 DX_L DX_R D_L D_R VDDHD VDDI VHI_VDD VLO_VDD VSSI WEB WEB3B X3B[0] 
+ X3B[1] X3B[2] X3B[3] X3B[4] X3B[5] X3B[6] X3B[7] X3B[8] X3B[9] X3B[10] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] Y3B[0] Y3B[1] Y3B[2] 
+ Y3B[3] Y[0] Y[1] Y[2] Y[3]
*.PININFO BWEB_L:I BWEB_R:I CEB:I CLK:I D_L:I D_R:I WEB:I X[0]:I X[1]:I X[2]:I 
*.PININFO X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I BWEBX_L:O BWEBX_R:O CEB3B:O CLK2:O DX_L:O 
*.PININFO DX_R:O VHI_VDD:O VLO_VDD:O WEB3B:O X3B[0]:O X3B[1]:O X3B[2]:O 
*.PININFO X3B[3]:O X3B[4]:O X3B[5]:O X3B[6]:O X3B[7]:O X3B[8]:O X3B[9]:O 
*.PININFO X3B[10]:O Y3B[0]:O Y3B[1]:O Y3B[2]:O Y3B[3]:O VDDHD:B VDDI:B VSSI:B
XBIST_CEB CEB CEB3B VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_WEB WEB WEB3B VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[0] X[0] X3B[0] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[1] X[1] X3B[1] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[2] X[2] X3B[2] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[3] X[3] X3B[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[4] X[4] X3B[4] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[5] X[5] X3B[5] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[6] X[6] X3B[6] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[7] X[7] X3B[7] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[8] X[8] X3B[8] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[9] X[9] X3B[9] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_X[10] X[10] X3B[10] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_Y[0] Y[0] Y3B[0] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_Y[1] Y[1] Y3B[1] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_Y[2] Y[2] Y3B[2] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XBIST_Y[3] Y[3] Y3B[3] VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST
XVHILO VDDI VHI_VDD VLO_VDD VSSI S1BSVTSWSO8000Y24_BIST_VHILO_M8_WOWO
XCLK_BUF CLK CLK2 VDDHD VDDI VSSI S1BSVTSWSO8000Y24_CLK_BUF
XIO_BIST_L_L BWEB_L BWEBX_L D_L DX_L VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST_WOLS_IO
XIO_BIST_LS_R BWEB_R BWEBX_R D_R DX_R VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST_WOLS_IO
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    CNT_M16_IOX2_WOBIST_SR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_CNT_M16_IOX2_WOBIST_SR AWT AWT2 BLTRKWLDRV BWEB_L BWEB_R CEB CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DSLP_BUF D_L D_R GBLB_L GBLB_R GBL_L GBL_R GWB_L GWB_R GW_L GW_R Q_L Q_R RE 
+ RTSEL[0] RTSEL[1] SD SLP SLP_BUF SLP_LBACK SLP_LCTRL SLP_Q SLP_RBACK TK TM 
+ TRKBL VDDHD VDDI VHI VHI_VDD VLO VLO_VDD VSSI WE WEB WLP_SAE WLP_SAEB 
+ WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] 
+ X[7] X[8] X[9] X[10] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1]
*.PININFO AWT:I BWEB_L:I BWEB_R:I CEB:I CLK:I D_L:I D_R:I GBLB_L:I GBLB_R:I 
*.PININFO GBL_L:I GBL_R:I RTSEL[0]:I RTSEL[1]:I SD:I SLP:I TM:I WEB:I 
*.PININFO WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I 
*.PININFO X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I Y[0]:I Y[1]:I Y[2]:I 
*.PININFO Y[3]:I AWT2:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O 
*.PININFO DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O 
*.PININFO DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O 
*.PININFO DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O 
*.PININFO DEC_X2[2]:O DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O 
*.PININFO DEC_X3[3]:O DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O 
*.PININFO DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O 
*.PININFO DEC_Y[6]:O DEC_Y[7]:O DSLP_BUF:O GWB_L:O GWB_R:O GW_L:O GW_R:O Q_L:O 
*.PININFO Q_R:O RE:O SLP_BUF:O SLP_LCTRL:O SLP_Q:O TK:O TRKBL:O WE:O WLP_SAE:O 
*.PININFO WLP_SAEB:O WLP_SAE_TK:O YL[0]:O YL[1]:O SLP_LBACK:B SLP_RBACK:B 
*.PININFO VDDHD:B VDDI:B VHI:B VHI_VDD:B VLO:B VLO_VDD:B VSSI:B
XCNTIO AWT AWT2 BLTRKWLDRV NET0108 NET084 BWEBX_L BWEBX_R CEB3B NET088 CKD 
+ CLK2 CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] 
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] 
+ DEC_Y[7] NET239 NET0116 NET253 DSLP_BUF DX_L DX_R GBLB_L GBLB_R GBL_L GBL_R 
+ GWB_L GWB_R GW_L GW_R NET249 Q_L Q_R RE NET0120 NET0100 RTSEL[0] RTSEL[1] SD 
+ NET063 SLP SLP_BUF SLP_LBACK SLP_LCTRL SLP_Q SLP_RBACK TK TM TRKBL VDDI 
+ VDDHD VDDHD VDDI VHI VLO VSSI WE WEB3B NET0106 WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] X3B[0] X3B[1] X3B[2] X3B[3] X3B[4] X3B[5] X3B[6] 
+ X3B[7] X3B[8] X3B[9] X3B[10] NET252 NET252 NET252 NET252 NET252 NET252 
+ NET252 NET252 NET252 NET252 NET252 Y3B[0] Y3B[1] Y3B[2] Y3B[3] YL[0] YL[1] 
+ NET246 NET246 NET246 NET246 S1BSVTSWSO8000Y24_CNT_M16_IOX2_WOBIST
XCNT_BIST_LS BWEBX_L BWEBX_R BWEB_L BWEB_R CEB CEB3B CLK CLK2 DX_L DX_R D_L 
+ D_R VDDHD VDDI VHI_VDD VLO_VDD VSSI WEB WEB3B X3B[0] X3B[1] X3B[2] X3B[3] 
+ X3B[4] X3B[5] X3B[6] X3B[7] X3B[8] X3B[9] X3B[10] X[0] X[1] X[2] X[3] X[4] 
+ X[5] X[6] X[7] X[8] X[9] X[10] Y3B[0] Y3B[1] Y3B[2] Y3B[3] Y[0] Y[1] Y[2] 
+ Y[3] S1BSVTSWSO8000Y24_WOBIST_WOLS_CNT_M16_IOX2
.ENDS

************************************************************************
* LIBRARY NAME: N28HP_SP_LEAFCELLS
* CELL NAME:    IO_M16_WOBIST_SR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1BSVTSWSO8000Y24_IO_M16_WOBIST_SR AWT BWEB CKD D GBL GBLB GW GWB IOPD PDI PDO Q SLP_Q 
+ VDDHD VDDI VSSI WLP_SAEB
*.PININFO AWT:I BWEB:I CKD:I D:I SLP_Q:I WLP_SAEB:I GW:O GWB:O PDO:O Q:O GBL:B 
*.PININFO GBLB:B IOPD:B PDI:B VDDHD:B VDDI:B VSSI:B
XI163 AWT BWEBX NET025 CKD DX NET026 GBL GBLB GW GWB IOPD PDI PDO Q SLP_Q VDDI 
+ VDDHD VDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16_WOBIST
XWOBIST_WOLS_IO BWEB BWEBX D DX VDDHD VDDI VSSI S1BSVTSWSO8000Y24_WOBIST_WOLS_IO
.ENDS




**** End of leaf cells

.SUBCKT S1BSVTSWSO8000Y24_CELL_ARR_X BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6]
+ BL[7] BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17]
+ BL[18] BL[19] BL[20] BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28]
+ BL[29] BL[30] BL[31] BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39]
+ BL[40] BL[41] BL[42] BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50]
+ BL[51] BL[52] BL[53] BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61]
+ BL[62] BL[63] BL[64] BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72]
+ BL[73] BL[74] BL[75] BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83]
+ BL[84] BL[85] BL[86] BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94]
+ BL[95] BL[96] BL[97] BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104]
+ BL[105] BL[106] BL[107] BL[108] BL[109] BL[110] BL[111] BL[112] BL[113]
+ BL[114] BL[115] BL[116] BL[117] BL[118] BL[119] BL[120] BL[121] BL[122]
+ BL[123] BL[124] BL[125] BL[126] BL[127] BL[128] BL[129] BL[130] BL[131]
+ BL[132] BL[133] BL[134] BL[135] BL[136] BL[137] BL[138] BL[139] BL[140]
+ BL[141] BL[142] BL[143] BL[144] BL[145] BL[146] BL[147] BL[148] BL[149]
+ BL[150] BL[151] BL[152] BL[153] BL[154] BL[155] BL[156] BL[157] BL[158]
+ BL[159] BL[160] BL[161] BL[162] BL[163] BL[164] BL[165] BL[166] BL[167]
+ BL[168] BL[169] BL[170] BL[171] BL[172] BL[173] BL[174] BL[175] BL[176]
+ BL[177] BL[178] BL[179] BL[180] BL[181] BL[182] BL[183] BL[184] BL[185]
+ BL[186] BL[187] BL[188] BL[189] BL[190] BL[191] BL[192] BL[193] BL[194]
+ BL[195] BL[196] BL[197] BL[198] BL[199] BL[200] BL[201] BL[202] BL[203]
+ BL[204] BL[205] BL[206] BL[207] BL[208] BL[209] BL[210] BL[211] BL[212]
+ BL[213] BL[214] BL[215] BL[216] BL[217] BL[218] BL[219] BL[220] BL[221]
+ BL[222] BL[223] BL[224] BL[225] BL[226] BL[227] BL[228] BL[229] BL[230]
+ BL[231] BL[232] BL[233] BL[234] BL[235] BL[236] BL[237] BL[238] BL[239]
+ BL[240] BL[241] BL[242] BL[243] BL[244] BL[245] BL[246] BL[247] BL[248]
+ BL[249] BL[250] BL[251] BL[252] BL[253] BL[254] BL[255] BL[256] BL[257]
+ BL[258] BL[259] BL[260] BL[261] BL[262] BL[263] BL[264] BL[265] BL[266]
+ BL[267] BL[268] BL[269] BL[270] BL[271] BL[272] BL[273] BL[274] BL[275]
+ BL[276] BL[277] BL[278] BL[279] BL[280] BL[281] BL[282] BL[283] BL[284]
+ BL[285] BL[286] BL[287] BL[288] BL[289] BL[290] BL[291] BL[292] BL[293]
+ BL[294] BL[295] BL[296] BL[297] BL[298] BL[299] BL[300] BL[301] BL[302]
+ BL[303] BL[304] BL[305] BL[306] BL[307] BL[308] BL[309] BL[310] BL[311]
+ BL[312] BL[313] BL[314] BL[315] BL[316] BL[317] BL[318] BL[319] BL[320]
+ BL[321] BL[322] BL[323] BL[324] BL[325] BL[326] BL[327] BL[328] BL[329]
+ BL[330] BL[331] BL[332] BL[333] BL[334] BL[335] BL[336] BL[337] BL[338]
+ BL[339] BL[340] BL[341] BL[342] BL[343] BL[344] BL[345] BL[346] BL[347]
+ BL[348] BL[349] BL[350] BL[351] BL[352] BL[353] BL[354] BL[355] BL[356]
+ BL[357] BL[358] BL[359] BL[360] BL[361] BL[362] BL[363] BL[364] BL[365]
+ BL[366] BL[367] BL[368] BL[369] BL[370] BL[371] BL[372] BL[373] BL[374]
+ BL[375] BL[376] BL[377] BL[378] BL[379] BL[380] BL[381] BL[382] BL[383]
+ BL[384] BL[385] BL[386] BL[387] BL[388] BL[389] BL[390] BL[391] BL[392]
+ BL[393] BL[394] BL[395] BL[396] BL[397] BL[398] BL[399] BL[400] BL[401]
+ BL[402] BL[403] BL[404] BL[405] BL[406] BL[407] BL[408] BL[409] BL[410]
+ BL[411] BL[412] BL[413] BL[414] BL[415] BL[416] BL[417] BL[418] BL[419]
+ BL[420] BL[421] BL[422] BL[423] BL[424] BL[425] BL[426] BL[427] BL[428]
+ BL[429] BL[430] BL[431] BL[432] BL[433] BL[434] BL[435] BL[436] BL[437]
+ BL[438] BL[439] BL[440] BL[441] BL[442] BL[443] BL[444] BL[445] BL[446]
+ BL[447] BL[448] BL[449] BL[450] BL[451] BL[452] BL[453] BL[454] BL[455]
+ BL[456] BL[457] BL[458] BL[459] BL[460] BL[461] BL[462] BL[463] BL[464]
+ BL[465] BL[466] BL[467] BL[468] BL[469] BL[470] BL[471] BL[472] BL[473]
+ BL[474] BL[475] BL[476] BL[477] BL[478] BL[479] BL[480] BL[481] BL[482]
+ BL[483] BL[484] BL[485] BL[486] BL[487] BL[488] BL[489] BL[490] BL[491]
+ BL[492] BL[493] BL[494] BL[495] BL[496] BL[497] BL[498] BL[499] BL[500]
+ BL[501] BL[502] BL[503] BL[504] BL[505] BL[506] BL[507] BL[508] BL[509]
+ BL[510] BL[511] BL[512] BL[513] BL[514] BL[515] BL[516] BL[517] BL[518]
+ BL[519] BL[520] BL[521] BL[522] BL[523] BL[524] BL[525] BL[526] BL[527]
+ BL[528] BL[529] BL[530] BL[531] BL[532] BL[533] BL[534] BL[535] BL[536]
+ BL[537] BL[538] BL[539] BL[540] BL[541] BL[542] BL[543] BL[544] BL[545]
+ BL[546] BL[547] BL[548] BL[549] BL[550] BL[551] BL[552] BL[553] BL[554]
+ BL[555] BL[556] BL[557] BL[558] BL[559] BL[560] BL[561] BL[562] BL[563]
+ BL[564] BL[565] BL[566] BL[567] BL[568] BL[569] BL[570] BL[571] BL[572]
+ BL[573] BL[574] BL[575] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] BLB[256] BLB[257] BLB[258]
+ BLB[259] BLB[260] BLB[261] BLB[262] BLB[263] BLB[264] BLB[265] BLB[266]
+ BLB[267] BLB[268] BLB[269] BLB[270] BLB[271] BLB[272] BLB[273] BLB[274]
+ BLB[275] BLB[276] BLB[277] BLB[278] BLB[279] BLB[280] BLB[281] BLB[282]
+ BLB[283] BLB[284] BLB[285] BLB[286] BLB[287] BLB[288] BLB[289] BLB[290]
+ BLB[291] BLB[292] BLB[293] BLB[294] BLB[295] BLB[296] BLB[297] BLB[298]
+ BLB[299] BLB[300] BLB[301] BLB[302] BLB[303] BLB[304] BLB[305] BLB[306]
+ BLB[307] BLB[308] BLB[309] BLB[310] BLB[311] BLB[312] BLB[313] BLB[314]
+ BLB[315] BLB[316] BLB[317] BLB[318] BLB[319] BLB[320] BLB[321] BLB[322]
+ BLB[323] BLB[324] BLB[325] BLB[326] BLB[327] BLB[328] BLB[329] BLB[330]
+ BLB[331] BLB[332] BLB[333] BLB[334] BLB[335] BLB[336] BLB[337] BLB[338]
+ BLB[339] BLB[340] BLB[341] BLB[342] BLB[343] BLB[344] BLB[345] BLB[346]
+ BLB[347] BLB[348] BLB[349] BLB[350] BLB[351] BLB[352] BLB[353] BLB[354]
+ BLB[355] BLB[356] BLB[357] BLB[358] BLB[359] BLB[360] BLB[361] BLB[362]
+ BLB[363] BLB[364] BLB[365] BLB[366] BLB[367] BLB[368] BLB[369] BLB[370]
+ BLB[371] BLB[372] BLB[373] BLB[374] BLB[375] BLB[376] BLB[377] BLB[378]
+ BLB[379] BLB[380] BLB[381] BLB[382] BLB[383] BLB[384] BLB[385] BLB[386]
+ BLB[387] BLB[388] BLB[389] BLB[390] BLB[391] BLB[392] BLB[393] BLB[394]
+ BLB[395] BLB[396] BLB[397] BLB[398] BLB[399] BLB[400] BLB[401] BLB[402]
+ BLB[403] BLB[404] BLB[405] BLB[406] BLB[407] BLB[408] BLB[409] BLB[410]
+ BLB[411] BLB[412] BLB[413] BLB[414] BLB[415] BLB[416] BLB[417] BLB[418]
+ BLB[419] BLB[420] BLB[421] BLB[422] BLB[423] BLB[424] BLB[425] BLB[426]
+ BLB[427] BLB[428] BLB[429] BLB[430] BLB[431] BLB[432] BLB[433] BLB[434]
+ BLB[435] BLB[436] BLB[437] BLB[438] BLB[439] BLB[440] BLB[441] BLB[442]
+ BLB[443] BLB[444] BLB[445] BLB[446] BLB[447] BLB[448] BLB[449] BLB[450]
+ BLB[451] BLB[452] BLB[453] BLB[454] BLB[455] BLB[456] BLB[457] BLB[458]
+ BLB[459] BLB[460] BLB[461] BLB[462] BLB[463] BLB[464] BLB[465] BLB[466]
+ BLB[467] BLB[468] BLB[469] BLB[470] BLB[471] BLB[472] BLB[473] BLB[474]
+ BLB[475] BLB[476] BLB[477] BLB[478] BLB[479] BLB[480] BLB[481] BLB[482]
+ BLB[483] BLB[484] BLB[485] BLB[486] BLB[487] BLB[488] BLB[489] BLB[490]
+ BLB[491] BLB[492] BLB[493] BLB[494] BLB[495] BLB[496] BLB[497] BLB[498]
+ BLB[499] BLB[500] BLB[501] BLB[502] BLB[503] BLB[504] BLB[505] BLB[506]
+ BLB[507] BLB[508] BLB[509] BLB[510] BLB[511] BLB[512] BLB[513] BLB[514]
+ BLB[515] BLB[516] BLB[517] BLB[518] BLB[519] BLB[520] BLB[521] BLB[522]
+ BLB[523] BLB[524] BLB[525] BLB[526] BLB[527] BLB[528] BLB[529] BLB[530]
+ BLB[531] BLB[532] BLB[533] BLB[534] BLB[535] BLB[536] BLB[537] BLB[538]
+ BLB[539] BLB[540] BLB[541] BLB[542] BLB[543] BLB[544] BLB[545] BLB[546]
+ BLB[547] BLB[548] BLB[549] BLB[550] BLB[551] BLB[552] BLB[553] BLB[554]
+ BLB[555] BLB[556] BLB[557] BLB[558] BLB[559] BLB[560] BLB[561] BLB[562]
+ BLB[563] BLB[564] BLB[565] BLB[566] BLB[567] BLB[568] BLB[569] BLB[570]
+ BLB[571] BLB[572] BLB[573] BLB[574] BLB[575] WL[0] WL[1] VXDDAI VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10]
+ GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21]
+ GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32]
+ GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
XMCB_0 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10] BL[11]
+ BL[12] BL[13] BL[14] BL[15] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] GBL[0]
+ GBLB[0] GW[0] GWB[0] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_1 BL[16] BL[17] BL[18] BL[19] BL[20] BL[21] BL[22] BL[23] BL[24] BL[25]
+ BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BLB[16] BLB[17] BLB[18] BLB[19]
+ BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28]
+ BLB[29] BLB[30] BLB[31] GBL[1] GBLB[1] GW[1] GWB[1] VXDDAI VDDI VSSI WL[0]
+ WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_2 BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41]
+ BL[42] BL[43] BL[44] BL[45] BL[46] BL[47] BLB[32] BLB[33] BLB[34] BLB[35]
+ BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44]
+ BLB[45] BLB[46] BLB[47] GBL[2] GBLB[2] GW[2] GWB[2] VXDDAI VDDI VSSI WL[0]
+ WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_3 BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54] BL[55] BL[56] BL[57]
+ BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] GBL[3] GBLB[3] GW[3] GWB[3] VXDDAI VDDI VSSI WL[0]
+ WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_4 BL[64] BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73]
+ BL[74] BL[75] BL[76] BL[77] BL[78] BL[79] BLB[64] BLB[65] BLB[66] BLB[67]
+ BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76]
+ BLB[77] BLB[78] BLB[79] GBL[4] GBLB[4] GW[4] GWB[4] VXDDAI VDDI VSSI WL[0]
+ WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_5 BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87] BL[88] BL[89]
+ BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] GBL[5] GBLB[5] GW[5] GWB[5] VXDDAI VDDI VSSI WL[0]
+ WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_6 BL[96] BL[97] BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104]
+ BL[105] BL[106] BL[107] BL[108] BL[109] BL[110] BL[111] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] GBL[6] GBLB[6] GW[6] GWB[6]
+ VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_7 BL[112] BL[113] BL[114] BL[115] BL[116] BL[117] BL[118] BL[119] BL[120]
+ BL[121] BL[122] BL[123] BL[124] BL[125] BL[126] BL[127] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] GBL[7] GBLB[7] GW[7]
+ GWB[7] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_8 BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135] BL[136]
+ BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] GBL[8] GBLB[8] GW[8]
+ GWB[8] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_9 BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] GBL[9] GBLB[9] GW[9]
+ GWB[9] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_10 BL[160] BL[161] BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168]
+ BL[169] BL[170] BL[171] BL[172] BL[173] BL[174] BL[175] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] GBL[10] GBLB[10] GW[10]
+ GWB[10] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_11 BL[176] BL[177] BL[178] BL[179] BL[180] BL[181] BL[182] BL[183] BL[184]
+ BL[185] BL[186] BL[187] BL[188] BL[189] BL[190] BL[191] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] GBL[11] GBLB[11] GW[11]
+ GWB[11] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_12 BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198] BL[199] BL[200]
+ BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] GBL[12] GBLB[12] GW[12]
+ GWB[12] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_13 BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] GBL[13] GBLB[13] GW[13]
+ GWB[13] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_14 BL[224] BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232]
+ BL[233] BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] GBL[14] GBLB[14] GW[14]
+ GWB[14] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_15 BL[240] BL[241] BL[242] BL[243] BL[244] BL[245] BL[246] BL[247] BL[248]
+ BL[249] BL[250] BL[251] BL[252] BL[253] BL[254] BL[255] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] GBL[15] GBLB[15] GW[15]
+ GWB[15] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_16 BL[256] BL[257] BL[258] BL[259] BL[260] BL[261] BL[262] BL[263] BL[264]
+ BL[265] BL[266] BL[267] BL[268] BL[269] BL[270] BL[271] BLB[256] BLB[257]
+ BLB[258] BLB[259] BLB[260] BLB[261] BLB[262] BLB[263] BLB[264] BLB[265]
+ BLB[266] BLB[267] BLB[268] BLB[269] BLB[270] BLB[271] GBL[16] GBLB[16] GW[16]
+ GWB[16] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_17 BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279] BL[280]
+ BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BLB[272] BLB[273]
+ BLB[274] BLB[275] BLB[276] BLB[277] BLB[278] BLB[279] BLB[280] BLB[281]
+ BLB[282] BLB[283] BLB[284] BLB[285] BLB[286] BLB[287] GBL[17] GBLB[17] GW[17]
+ GWB[17] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_18 BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BLB[288] BLB[289]
+ BLB[290] BLB[291] BLB[292] BLB[293] BLB[294] BLB[295] BLB[296] BLB[297]
+ BLB[298] BLB[299] BLB[300] BLB[301] BLB[302] BLB[303] GBL[18] GBLB[18] GW[18]
+ GWB[18] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_19 BL[304] BL[305] BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312]
+ BL[313] BL[314] BL[315] BL[316] BL[317] BL[318] BL[319] BLB[304] BLB[305]
+ BLB[306] BLB[307] BLB[308] BLB[309] BLB[310] BLB[311] BLB[312] BLB[313]
+ BLB[314] BLB[315] BLB[316] BLB[317] BLB[318] BLB[319] GBL[19] GBLB[19] GW[19]
+ GWB[19] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_20 BL[320] BL[321] BL[322] BL[323] BL[324] BL[325] BL[326] BL[327] BL[328]
+ BL[329] BL[330] BL[331] BL[332] BL[333] BL[334] BL[335] BLB[320] BLB[321]
+ BLB[322] BLB[323] BLB[324] BLB[325] BLB[326] BLB[327] BLB[328] BLB[329]
+ BLB[330] BLB[331] BLB[332] BLB[333] BLB[334] BLB[335] GBL[20] GBLB[20] GW[20]
+ GWB[20] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_21 BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342] BL[343] BL[344]
+ BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351] BLB[336] BLB[337]
+ BLB[338] BLB[339] BLB[340] BLB[341] BLB[342] BLB[343] BLB[344] BLB[345]
+ BLB[346] BLB[347] BLB[348] BLB[349] BLB[350] BLB[351] GBL[21] GBLB[21] GW[21]
+ GWB[21] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_22 BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BLB[352] BLB[353]
+ BLB[354] BLB[355] BLB[356] BLB[357] BLB[358] BLB[359] BLB[360] BLB[361]
+ BLB[362] BLB[363] BLB[364] BLB[365] BLB[366] BLB[367] GBL[22] GBLB[22] GW[22]
+ GWB[22] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_23 BL[368] BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376]
+ BL[377] BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BLB[368] BLB[369]
+ BLB[370] BLB[371] BLB[372] BLB[373] BLB[374] BLB[375] BLB[376] BLB[377]
+ BLB[378] BLB[379] BLB[380] BLB[381] BLB[382] BLB[383] GBL[23] GBLB[23] GW[23]
+ GWB[23] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_24 BL[384] BL[385] BL[386] BL[387] BL[388] BL[389] BL[390] BL[391] BL[392]
+ BL[393] BL[394] BL[395] BL[396] BL[397] BL[398] BL[399] BLB[384] BLB[385]
+ BLB[386] BLB[387] BLB[388] BLB[389] BLB[390] BLB[391] BLB[392] BLB[393]
+ BLB[394] BLB[395] BLB[396] BLB[397] BLB[398] BLB[399] GBL[24] GBLB[24] GW[24]
+ GWB[24] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_25 BL[400] BL[401] BL[402] BL[403] BL[404] BL[405] BL[406] BL[407] BL[408]
+ BL[409] BL[410] BL[411] BL[412] BL[413] BL[414] BL[415] BLB[400] BLB[401]
+ BLB[402] BLB[403] BLB[404] BLB[405] BLB[406] BLB[407] BLB[408] BLB[409]
+ BLB[410] BLB[411] BLB[412] BLB[413] BLB[414] BLB[415] GBL[25] GBLB[25] GW[25]
+ GWB[25] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_26 BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423] BL[424]
+ BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BLB[416] BLB[417]
+ BLB[418] BLB[419] BLB[420] BLB[421] BLB[422] BLB[423] BLB[424] BLB[425]
+ BLB[426] BLB[427] BLB[428] BLB[429] BLB[430] BLB[431] GBL[26] GBLB[26] GW[26]
+ GWB[26] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_27 BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BLB[432] BLB[433]
+ BLB[434] BLB[435] BLB[436] BLB[437] BLB[438] BLB[439] BLB[440] BLB[441]
+ BLB[442] BLB[443] BLB[444] BLB[445] BLB[446] BLB[447] GBL[27] GBLB[27] GW[27]
+ GWB[27] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_28 BL[448] BL[449] BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456]
+ BL[457] BL[458] BL[459] BL[460] BL[461] BL[462] BL[463] BLB[448] BLB[449]
+ BLB[450] BLB[451] BLB[452] BLB[453] BLB[454] BLB[455] BLB[456] BLB[457]
+ BLB[458] BLB[459] BLB[460] BLB[461] BLB[462] BLB[463] GBL[28] GBLB[28] GW[28]
+ GWB[28] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_29 BL[464] BL[465] BL[466] BL[467] BL[468] BL[469] BL[470] BL[471] BL[472]
+ BL[473] BL[474] BL[475] BL[476] BL[477] BL[478] BL[479] BLB[464] BLB[465]
+ BLB[466] BLB[467] BLB[468] BLB[469] BLB[470] BLB[471] BLB[472] BLB[473]
+ BLB[474] BLB[475] BLB[476] BLB[477] BLB[478] BLB[479] GBL[29] GBLB[29] GW[29]
+ GWB[29] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_30 BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486] BL[487] BL[488]
+ BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495] BLB[480] BLB[481]
+ BLB[482] BLB[483] BLB[484] BLB[485] BLB[486] BLB[487] BLB[488] BLB[489]
+ BLB[490] BLB[491] BLB[492] BLB[493] BLB[494] BLB[495] GBL[30] GBLB[30] GW[30]
+ GWB[30] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_31 BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BLB[496] BLB[497]
+ BLB[498] BLB[499] BLB[500] BLB[501] BLB[502] BLB[503] BLB[504] BLB[505]
+ BLB[506] BLB[507] BLB[508] BLB[509] BLB[510] BLB[511] GBL[31] GBLB[31] GW[31]
+ GWB[31] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_32 BL[512] BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520]
+ BL[521] BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BLB[512] BLB[513]
+ BLB[514] BLB[515] BLB[516] BLB[517] BLB[518] BLB[519] BLB[520] BLB[521]
+ BLB[522] BLB[523] BLB[524] BLB[525] BLB[526] BLB[527] GBL[32] GBLB[32] GW[32]
+ GWB[32] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_33 BL[528] BL[529] BL[530] BL[531] BL[532] BL[533] BL[534] BL[535] BL[536]
+ BL[537] BL[538] BL[539] BL[540] BL[541] BL[542] BL[543] BLB[528] BLB[529]
+ BLB[530] BLB[531] BLB[532] BLB[533] BLB[534] BLB[535] BLB[536] BLB[537]
+ BLB[538] BLB[539] BLB[540] BLB[541] BLB[542] BLB[543] GBL[33] GBLB[33] GW[33]
+ GWB[33] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_34 BL[544] BL[545] BL[546] BL[547] BL[548] BL[549] BL[550] BL[551] BL[552]
+ BL[553] BL[554] BL[555] BL[556] BL[557] BL[558] BL[559] BLB[544] BLB[545]
+ BLB[546] BLB[547] BLB[548] BLB[549] BLB[550] BLB[551] BLB[552] BLB[553]
+ BLB[554] BLB[555] BLB[556] BLB[557] BLB[558] BLB[559] GBL[34] GBLB[34] GW[34]
+ GWB[34] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
XMCB_35 BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567] BL[568]
+ BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[560] BLB[561]
+ BLB[562] BLB[563] BLB[564] BLB[565] BLB[566] BLB[567] BLB[568] BLB[569]
+ BLB[570] BLB[571] BLB[572] BLB[573] BLB[574] BLB[575] GBL[35] GBLB[35] GW[35]
+ GWB[35] VXDDAI VDDI VSSI WL[0] WL[1] S1BSVTSWSO8000Y24_MCB_2X16
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_CELL_ARR_XY_F BL[0] BL[1] BL[2] BL[3] BL[4] BL[5]
+ BL[6] BL[7] BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16]
+ BL[17] BL[18] BL[19] BL[20] BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27]
+ BL[28] BL[29] BL[30] BL[31] BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38]
+ BL[39] BL[40] BL[41] BL[42] BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49]
+ BL[50] BL[51] BL[52] BL[53] BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60]
+ BL[61] BL[62] BL[63] BL[64] BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71]
+ BL[72] BL[73] BL[74] BL[75] BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82]
+ BL[83] BL[84] BL[85] BL[86] BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93]
+ BL[94] BL[95] BL[96] BL[97] BL[98] BL[99] BL[100] BL[101] BL[102] BL[103]
+ BL[104] BL[105] BL[106] BL[107] BL[108] BL[109] BL[110] BL[111] BL[112]
+ BL[113] BL[114] BL[115] BL[116] BL[117] BL[118] BL[119] BL[120] BL[121]
+ BL[122] BL[123] BL[124] BL[125] BL[126] BL[127] BL[128] BL[129] BL[130]
+ BL[131] BL[132] BL[133] BL[134] BL[135] BL[136] BL[137] BL[138] BL[139]
+ BL[140] BL[141] BL[142] BL[143] BL[144] BL[145] BL[146] BL[147] BL[148]
+ BL[149] BL[150] BL[151] BL[152] BL[153] BL[154] BL[155] BL[156] BL[157]
+ BL[158] BL[159] BL[160] BL[161] BL[162] BL[163] BL[164] BL[165] BL[166]
+ BL[167] BL[168] BL[169] BL[170] BL[171] BL[172] BL[173] BL[174] BL[175]
+ BL[176] BL[177] BL[178] BL[179] BL[180] BL[181] BL[182] BL[183] BL[184]
+ BL[185] BL[186] BL[187] BL[188] BL[189] BL[190] BL[191] BL[192] BL[193]
+ BL[194] BL[195] BL[196] BL[197] BL[198] BL[199] BL[200] BL[201] BL[202]
+ BL[203] BL[204] BL[205] BL[206] BL[207] BL[208] BL[209] BL[210] BL[211]
+ BL[212] BL[213] BL[214] BL[215] BL[216] BL[217] BL[218] BL[219] BL[220]
+ BL[221] BL[222] BL[223] BL[224] BL[225] BL[226] BL[227] BL[228] BL[229]
+ BL[230] BL[231] BL[232] BL[233] BL[234] BL[235] BL[236] BL[237] BL[238]
+ BL[239] BL[240] BL[241] BL[242] BL[243] BL[244] BL[245] BL[246] BL[247]
+ BL[248] BL[249] BL[250] BL[251] BL[252] BL[253] BL[254] BL[255] BL[256]
+ BL[257] BL[258] BL[259] BL[260] BL[261] BL[262] BL[263] BL[264] BL[265]
+ BL[266] BL[267] BL[268] BL[269] BL[270] BL[271] BL[272] BL[273] BL[274]
+ BL[275] BL[276] BL[277] BL[278] BL[279] BL[280] BL[281] BL[282] BL[283]
+ BL[284] BL[285] BL[286] BL[287] BL[288] BL[289] BL[290] BL[291] BL[292]
+ BL[293] BL[294] BL[295] BL[296] BL[297] BL[298] BL[299] BL[300] BL[301]
+ BL[302] BL[303] BL[304] BL[305] BL[306] BL[307] BL[308] BL[309] BL[310]
+ BL[311] BL[312] BL[313] BL[314] BL[315] BL[316] BL[317] BL[318] BL[319]
+ BL[320] BL[321] BL[322] BL[323] BL[324] BL[325] BL[326] BL[327] BL[328]
+ BL[329] BL[330] BL[331] BL[332] BL[333] BL[334] BL[335] BL[336] BL[337]
+ BL[338] BL[339] BL[340] BL[341] BL[342] BL[343] BL[344] BL[345] BL[346]
+ BL[347] BL[348] BL[349] BL[350] BL[351] BL[352] BL[353] BL[354] BL[355]
+ BL[356] BL[357] BL[358] BL[359] BL[360] BL[361] BL[362] BL[363] BL[364]
+ BL[365] BL[366] BL[367] BL[368] BL[369] BL[370] BL[371] BL[372] BL[373]
+ BL[374] BL[375] BL[376] BL[377] BL[378] BL[379] BL[380] BL[381] BL[382]
+ BL[383] BL[384] BL[385] BL[386] BL[387] BL[388] BL[389] BL[390] BL[391]
+ BL[392] BL[393] BL[394] BL[395] BL[396] BL[397] BL[398] BL[399] BL[400]
+ BL[401] BL[402] BL[403] BL[404] BL[405] BL[406] BL[407] BL[408] BL[409]
+ BL[410] BL[411] BL[412] BL[413] BL[414] BL[415] BL[416] BL[417] BL[418]
+ BL[419] BL[420] BL[421] BL[422] BL[423] BL[424] BL[425] BL[426] BL[427]
+ BL[428] BL[429] BL[430] BL[431] BL[432] BL[433] BL[434] BL[435] BL[436]
+ BL[437] BL[438] BL[439] BL[440] BL[441] BL[442] BL[443] BL[444] BL[445]
+ BL[446] BL[447] BL[448] BL[449] BL[450] BL[451] BL[452] BL[453] BL[454]
+ BL[455] BL[456] BL[457] BL[458] BL[459] BL[460] BL[461] BL[462] BL[463]
+ BL[464] BL[465] BL[466] BL[467] BL[468] BL[469] BL[470] BL[471] BL[472]
+ BL[473] BL[474] BL[475] BL[476] BL[477] BL[478] BL[479] BL[480] BL[481]
+ BL[482] BL[483] BL[484] BL[485] BL[486] BL[487] BL[488] BL[489] BL[490]
+ BL[491] BL[492] BL[493] BL[494] BL[495] BL[496] BL[497] BL[498] BL[499]
+ BL[500] BL[501] BL[502] BL[503] BL[504] BL[505] BL[506] BL[507] BL[508]
+ BL[509] BL[510] BL[511] BL[512] BL[513] BL[514] BL[515] BL[516] BL[517]
+ BL[518] BL[519] BL[520] BL[521] BL[522] BL[523] BL[524] BL[525] BL[526]
+ BL[527] BL[528] BL[529] BL[530] BL[531] BL[532] BL[533] BL[534] BL[535]
+ BL[536] BL[537] BL[538] BL[539] BL[540] BL[541] BL[542] BL[543] BL[544]
+ BL[545] BL[546] BL[547] BL[548] BL[549] BL[550] BL[551] BL[552] BL[553]
+ BL[554] BL[555] BL[556] BL[557] BL[558] BL[559] BL[560] BL[561] BL[562]
+ BL[563] BL[564] BL[565] BL[566] BL[567] BL[568] BL[569] BL[570] BL[571]
+ BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] BLB[256] BLB[257]
+ BLB[258] BLB[259] BLB[260] BLB[261] BLB[262] BLB[263] BLB[264] BLB[265]
+ BLB[266] BLB[267] BLB[268] BLB[269] BLB[270] BLB[271] BLB[272] BLB[273]
+ BLB[274] BLB[275] BLB[276] BLB[277] BLB[278] BLB[279] BLB[280] BLB[281]
+ BLB[282] BLB[283] BLB[284] BLB[285] BLB[286] BLB[287] BLB[288] BLB[289]
+ BLB[290] BLB[291] BLB[292] BLB[293] BLB[294] BLB[295] BLB[296] BLB[297]
+ BLB[298] BLB[299] BLB[300] BLB[301] BLB[302] BLB[303] BLB[304] BLB[305]
+ BLB[306] BLB[307] BLB[308] BLB[309] BLB[310] BLB[311] BLB[312] BLB[313]
+ BLB[314] BLB[315] BLB[316] BLB[317] BLB[318] BLB[319] BLB[320] BLB[321]
+ BLB[322] BLB[323] BLB[324] BLB[325] BLB[326] BLB[327] BLB[328] BLB[329]
+ BLB[330] BLB[331] BLB[332] BLB[333] BLB[334] BLB[335] BLB[336] BLB[337]
+ BLB[338] BLB[339] BLB[340] BLB[341] BLB[342] BLB[343] BLB[344] BLB[345]
+ BLB[346] BLB[347] BLB[348] BLB[349] BLB[350] BLB[351] BLB[352] BLB[353]
+ BLB[354] BLB[355] BLB[356] BLB[357] BLB[358] BLB[359] BLB[360] BLB[361]
+ BLB[362] BLB[363] BLB[364] BLB[365] BLB[366] BLB[367] BLB[368] BLB[369]
+ BLB[370] BLB[371] BLB[372] BLB[373] BLB[374] BLB[375] BLB[376] BLB[377]
+ BLB[378] BLB[379] BLB[380] BLB[381] BLB[382] BLB[383] BLB[384] BLB[385]
+ BLB[386] BLB[387] BLB[388] BLB[389] BLB[390] BLB[391] BLB[392] BLB[393]
+ BLB[394] BLB[395] BLB[396] BLB[397] BLB[398] BLB[399] BLB[400] BLB[401]
+ BLB[402] BLB[403] BLB[404] BLB[405] BLB[406] BLB[407] BLB[408] BLB[409]
+ BLB[410] BLB[411] BLB[412] BLB[413] BLB[414] BLB[415] BLB[416] BLB[417]
+ BLB[418] BLB[419] BLB[420] BLB[421] BLB[422] BLB[423] BLB[424] BLB[425]
+ BLB[426] BLB[427] BLB[428] BLB[429] BLB[430] BLB[431] BLB[432] BLB[433]
+ BLB[434] BLB[435] BLB[436] BLB[437] BLB[438] BLB[439] BLB[440] BLB[441]
+ BLB[442] BLB[443] BLB[444] BLB[445] BLB[446] BLB[447] BLB[448] BLB[449]
+ BLB[450] BLB[451] BLB[452] BLB[453] BLB[454] BLB[455] BLB[456] BLB[457]
+ BLB[458] BLB[459] BLB[460] BLB[461] BLB[462] BLB[463] BLB[464] BLB[465]
+ BLB[466] BLB[467] BLB[468] BLB[469] BLB[470] BLB[471] BLB[472] BLB[473]
+ BLB[474] BLB[475] BLB[476] BLB[477] BLB[478] BLB[479] BLB[480] BLB[481]
+ BLB[482] BLB[483] BLB[484] BLB[485] BLB[486] BLB[487] BLB[488] BLB[489]
+ BLB[490] BLB[491] BLB[492] BLB[493] BLB[494] BLB[495] BLB[496] BLB[497]
+ BLB[498] BLB[499] BLB[500] BLB[501] BLB[502] BLB[503] BLB[504] BLB[505]
+ BLB[506] BLB[507] BLB[508] BLB[509] BLB[510] BLB[511] BLB[512] BLB[513]
+ BLB[514] BLB[515] BLB[516] BLB[517] BLB[518] BLB[519] BLB[520] BLB[521]
+ BLB[522] BLB[523] BLB[524] BLB[525] BLB[526] BLB[527] BLB[528] BLB[529]
+ BLB[530] BLB[531] BLB[532] BLB[533] BLB[534] BLB[535] BLB[536] BLB[537]
+ BLB[538] BLB[539] BLB[540] BLB[541] BLB[542] BLB[543] BLB[544] BLB[545]
+ BLB[546] BLB[547] BLB[548] BLB[549] BLB[550] BLB[551] BLB[552] BLB[553]
+ BLB[554] BLB[555] BLB[556] BLB[557] BLB[558] BLB[559] BLB[560] BLB[561]
+ BLB[562] BLB[563] BLB[564] BLB[565] BLB[566] BLB[567] BLB[568] BLB[569]
+ BLB[570] BLB[571] BLB[572] BLB[573] BLB[574] BLB[575] WL[0] WL[1] WL[2] WL[3]
+ WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15]
+ WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26]
+ WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37]
+ WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48]
+ WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59]
+ WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70]
+ WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81]
+ WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92]
+ WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102]
+ WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111]
+ WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120]
+ WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129]
+ WL[130] WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138]
+ WL[139] WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147]
+ WL[148] WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156]
+ WL[157] WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165]
+ WL[166] WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174]
+ WL[175] WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183]
+ WL[184] WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192]
+ WL[193] WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201]
+ WL[202] WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210]
+ WL[211] WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219]
+ WL[220] WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228]
+ WL[229] WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237]
+ WL[238] WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246]
+ WL[247] WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] VXDDAI
+ VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8]
+ GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9]
+ GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20]
+ GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31]
+ GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35]
XCELL_ARR_X_0 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512] BL[513]
+ BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521] BL[522]
+ BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530] BL[531]
+ BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539] BL[540]
+ BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548] BL[549]
+ BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557] BL[558]
+ BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567]
+ BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[0] WL[1] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_1 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512] BL[513]
+ BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521] BL[522]
+ BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530] BL[531]
+ BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539] BL[540]
+ BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548] BL[549]
+ BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557] BL[558]
+ BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567]
+ BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[2] WL[3] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_2 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512] BL[513]
+ BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521] BL[522]
+ BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530] BL[531]
+ BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539] BL[540]
+ BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548] BL[549]
+ BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557] BL[558]
+ BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567]
+ BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[4] WL[5] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_3 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512] BL[513]
+ BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521] BL[522]
+ BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530] BL[531]
+ BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539] BL[540]
+ BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548] BL[549]
+ BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557] BL[558]
+ BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567]
+ BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[6] WL[7] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_4 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512] BL[513]
+ BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521] BL[522]
+ BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530] BL[531]
+ BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539] BL[540]
+ BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548] BL[549]
+ BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557] BL[558]
+ BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567]
+ BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[8] WL[9] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_5 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512] BL[513]
+ BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521] BL[522]
+ BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530] BL[531]
+ BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539] BL[540]
+ BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548] BL[549]
+ BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557] BL[558]
+ BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567]
+ BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[10] WL[11] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_6 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512] BL[513]
+ BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521] BL[522]
+ BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530] BL[531]
+ BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539] BL[540]
+ BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548] BL[549]
+ BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557] BL[558]
+ BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567]
+ BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[12] WL[13] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_7 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512] BL[513]
+ BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521] BL[522]
+ BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530] BL[531]
+ BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539] BL[540]
+ BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548] BL[549]
+ BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557] BL[558]
+ BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567]
+ BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[14] WL[15] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_8 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512] BL[513]
+ BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521] BL[522]
+ BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530] BL[531]
+ BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539] BL[540]
+ BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548] BL[549]
+ BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557] BL[558]
+ BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567]
+ BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[16] WL[17] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_9 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260] BL[261]
+ BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269] BL[270]
+ BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278] BL[279]
+ BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287] BL[288]
+ BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296] BL[297]
+ BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305] BL[306]
+ BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314] BL[315]
+ BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323] BL[324]
+ BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332] BL[333]
+ BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341] BL[342]
+ BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350] BL[351]
+ BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359] BL[360]
+ BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368] BL[369]
+ BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377] BL[378]
+ BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386] BL[387]
+ BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395] BL[396]
+ BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404] BL[405]
+ BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413] BL[414]
+ BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422] BL[423]
+ BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431] BL[432]
+ BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440] BL[441]
+ BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449] BL[450]
+ BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458] BL[459]
+ BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467] BL[468]
+ BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476] BL[477]
+ BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485] BL[486]
+ BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494] BL[495]
+ BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503] BL[504]
+ BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512] BL[513]
+ BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521] BL[522]
+ BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530] BL[531]
+ BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539] BL[540]
+ BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548] BL[549]
+ BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557] BL[558]
+ BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566] BL[567]
+ BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0] BLB[1]
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[18] WL[19] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_10 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[20] WL[21] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_11 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[22] WL[23] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_12 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[24] WL[25] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_13 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[26] WL[27] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_14 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[28] WL[29] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_15 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[30] WL[31] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_16 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[32] WL[33] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_17 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[34] WL[35] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_18 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[36] WL[37] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_19 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[38] WL[39] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_20 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[40] WL[41] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_21 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[42] WL[43] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_22 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[44] WL[45] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_23 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[46] WL[47] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_24 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[48] WL[49] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_25 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[50] WL[51] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_26 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[52] WL[53] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_27 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[54] WL[55] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_28 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[56] WL[57] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_29 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[58] WL[59] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_30 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[60] WL[61] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_31 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[62] WL[63] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_32 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[64] WL[65] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_33 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[66] WL[67] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_34 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[68] WL[69] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_35 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[70] WL[71] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_36 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[72] WL[73] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_37 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[74] WL[75] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_38 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[76] WL[77] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_39 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[78] WL[79] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_40 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[80] WL[81] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_41 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[82] WL[83] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_42 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[84] WL[85] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_43 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[86] WL[87] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_44 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[88] WL[89] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_45 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[90] WL[91] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_46 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[92] WL[93] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_47 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[94] WL[95] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_48 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[96] WL[97] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_49 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[98] WL[99] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_50 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[100] WL[101] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_51 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[102] WL[103] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_52 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[104] WL[105] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_53 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[106] WL[107] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_54 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[108] WL[109] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_55 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[110] WL[111] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_56 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[112] WL[113] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_57 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[114] WL[115] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_58 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[116] WL[117] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_59 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[118] WL[119] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_60 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[120] WL[121] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_61 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[122] WL[123] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_62 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[124] WL[125] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_63 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[126] WL[127] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_64 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[128] WL[129] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_65 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[130] WL[131] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_66 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[132] WL[133] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_67 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[134] WL[135] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_68 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[136] WL[137] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_69 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[138] WL[139] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_70 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[140] WL[141] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_71 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[142] WL[143] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_72 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[144] WL[145] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_73 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[146] WL[147] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_74 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[148] WL[149] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_75 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[150] WL[151] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_76 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[152] WL[153] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_77 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[154] WL[155] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_78 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[156] WL[157] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_79 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[158] WL[159] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_80 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[160] WL[161] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_81 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[162] WL[163] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_82 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[164] WL[165] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_83 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[166] WL[167] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_84 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[168] WL[169] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_85 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[170] WL[171] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_86 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[172] WL[173] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_87 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[174] WL[175] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_88 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[176] WL[177] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_89 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[178] WL[179] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_90 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[180] WL[181] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_91 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[182] WL[183] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_92 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[184] WL[185] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_93 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[186] WL[187] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_94 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[188] WL[189] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_95 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[190] WL[191] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_96 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[192] WL[193] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_97 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[194] WL[195] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_98 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[196] WL[197] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_99 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[198] WL[199] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_100 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[200] WL[201] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_101 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[202] WL[203] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_102 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[204] WL[205] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_103 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[206] WL[207] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_104 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[208] WL[209] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_105 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[210] WL[211] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_106 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[212] WL[213] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_107 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[214] WL[215] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_108 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[216] WL[217] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_109 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[218] WL[219] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_110 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[220] WL[221] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_111 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[222] WL[223] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_112 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[224] WL[225] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_113 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[226] WL[227] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_114 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[228] WL[229] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_115 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[230] WL[231] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_116 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[232] WL[233] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_117 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[234] WL[235] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_118 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[236] WL[237] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_119 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[238] WL[239] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_120 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[240] WL[241] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_121 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[242] WL[243] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_122 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[244] WL[245] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_123 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[246] WL[247] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_124 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[248] WL[249] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_125 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[250] WL[251] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_126 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[252] WL[253] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
XCELL_ARR_X_127 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BL[256] BL[257] BL[258] BL[259] BL[260]
+ BL[261] BL[262] BL[263] BL[264] BL[265] BL[266] BL[267] BL[268] BL[269]
+ BL[270] BL[271] BL[272] BL[273] BL[274] BL[275] BL[276] BL[277] BL[278]
+ BL[279] BL[280] BL[281] BL[282] BL[283] BL[284] BL[285] BL[286] BL[287]
+ BL[288] BL[289] BL[290] BL[291] BL[292] BL[293] BL[294] BL[295] BL[296]
+ BL[297] BL[298] BL[299] BL[300] BL[301] BL[302] BL[303] BL[304] BL[305]
+ BL[306] BL[307] BL[308] BL[309] BL[310] BL[311] BL[312] BL[313] BL[314]
+ BL[315] BL[316] BL[317] BL[318] BL[319] BL[320] BL[321] BL[322] BL[323]
+ BL[324] BL[325] BL[326] BL[327] BL[328] BL[329] BL[330] BL[331] BL[332]
+ BL[333] BL[334] BL[335] BL[336] BL[337] BL[338] BL[339] BL[340] BL[341]
+ BL[342] BL[343] BL[344] BL[345] BL[346] BL[347] BL[348] BL[349] BL[350]
+ BL[351] BL[352] BL[353] BL[354] BL[355] BL[356] BL[357] BL[358] BL[359]
+ BL[360] BL[361] BL[362] BL[363] BL[364] BL[365] BL[366] BL[367] BL[368]
+ BL[369] BL[370] BL[371] BL[372] BL[373] BL[374] BL[375] BL[376] BL[377]
+ BL[378] BL[379] BL[380] BL[381] BL[382] BL[383] BL[384] BL[385] BL[386]
+ BL[387] BL[388] BL[389] BL[390] BL[391] BL[392] BL[393] BL[394] BL[395]
+ BL[396] BL[397] BL[398] BL[399] BL[400] BL[401] BL[402] BL[403] BL[404]
+ BL[405] BL[406] BL[407] BL[408] BL[409] BL[410] BL[411] BL[412] BL[413]
+ BL[414] BL[415] BL[416] BL[417] BL[418] BL[419] BL[420] BL[421] BL[422]
+ BL[423] BL[424] BL[425] BL[426] BL[427] BL[428] BL[429] BL[430] BL[431]
+ BL[432] BL[433] BL[434] BL[435] BL[436] BL[437] BL[438] BL[439] BL[440]
+ BL[441] BL[442] BL[443] BL[444] BL[445] BL[446] BL[447] BL[448] BL[449]
+ BL[450] BL[451] BL[452] BL[453] BL[454] BL[455] BL[456] BL[457] BL[458]
+ BL[459] BL[460] BL[461] BL[462] BL[463] BL[464] BL[465] BL[466] BL[467]
+ BL[468] BL[469] BL[470] BL[471] BL[472] BL[473] BL[474] BL[475] BL[476]
+ BL[477] BL[478] BL[479] BL[480] BL[481] BL[482] BL[483] BL[484] BL[485]
+ BL[486] BL[487] BL[488] BL[489] BL[490] BL[491] BL[492] BL[493] BL[494]
+ BL[495] BL[496] BL[497] BL[498] BL[499] BL[500] BL[501] BL[502] BL[503]
+ BL[504] BL[505] BL[506] BL[507] BL[508] BL[509] BL[510] BL[511] BL[512]
+ BL[513] BL[514] BL[515] BL[516] BL[517] BL[518] BL[519] BL[520] BL[521]
+ BL[522] BL[523] BL[524] BL[525] BL[526] BL[527] BL[528] BL[529] BL[530]
+ BL[531] BL[532] BL[533] BL[534] BL[535] BL[536] BL[537] BL[538] BL[539]
+ BL[540] BL[541] BL[542] BL[543] BL[544] BL[545] BL[546] BL[547] BL[548]
+ BL[549] BL[550] BL[551] BL[552] BL[553] BL[554] BL[555] BL[556] BL[557]
+ BL[558] BL[559] BL[560] BL[561] BL[562] BL[563] BL[564] BL[565] BL[566]
+ BL[567] BL[568] BL[569] BL[570] BL[571] BL[572] BL[573] BL[574] BL[575] BLB[0]
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11]
+ BLB[12] BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20]
+ BLB[21] BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29]
+ BLB[30] BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38]
+ BLB[39] BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47]
+ BLB[48] BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56]
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65]
+ BLB[66] BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74]
+ BLB[75] BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83]
+ BLB[84] BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92]
+ BLB[93] BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101]
+ BLB[102] BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109]
+ BLB[110] BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117]
+ BLB[118] BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125]
+ BLB[126] BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133]
+ BLB[134] BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141]
+ BLB[142] BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149]
+ BLB[150] BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157]
+ BLB[158] BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165]
+ BLB[166] BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173]
+ BLB[174] BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181]
+ BLB[182] BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189]
+ BLB[190] BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197]
+ BLB[198] BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205]
+ BLB[206] BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213]
+ BLB[214] BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221]
+ BLB[222] BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229]
+ BLB[230] BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237]
+ BLB[238] BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245]
+ BLB[246] BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253]
+ BLB[254] BLB[255] BLB[256] BLB[257] BLB[258] BLB[259] BLB[260] BLB[261]
+ BLB[262] BLB[263] BLB[264] BLB[265] BLB[266] BLB[267] BLB[268] BLB[269]
+ BLB[270] BLB[271] BLB[272] BLB[273] BLB[274] BLB[275] BLB[276] BLB[277]
+ BLB[278] BLB[279] BLB[280] BLB[281] BLB[282] BLB[283] BLB[284] BLB[285]
+ BLB[286] BLB[287] BLB[288] BLB[289] BLB[290] BLB[291] BLB[292] BLB[293]
+ BLB[294] BLB[295] BLB[296] BLB[297] BLB[298] BLB[299] BLB[300] BLB[301]
+ BLB[302] BLB[303] BLB[304] BLB[305] BLB[306] BLB[307] BLB[308] BLB[309]
+ BLB[310] BLB[311] BLB[312] BLB[313] BLB[314] BLB[315] BLB[316] BLB[317]
+ BLB[318] BLB[319] BLB[320] BLB[321] BLB[322] BLB[323] BLB[324] BLB[325]
+ BLB[326] BLB[327] BLB[328] BLB[329] BLB[330] BLB[331] BLB[332] BLB[333]
+ BLB[334] BLB[335] BLB[336] BLB[337] BLB[338] BLB[339] BLB[340] BLB[341]
+ BLB[342] BLB[343] BLB[344] BLB[345] BLB[346] BLB[347] BLB[348] BLB[349]
+ BLB[350] BLB[351] BLB[352] BLB[353] BLB[354] BLB[355] BLB[356] BLB[357]
+ BLB[358] BLB[359] BLB[360] BLB[361] BLB[362] BLB[363] BLB[364] BLB[365]
+ BLB[366] BLB[367] BLB[368] BLB[369] BLB[370] BLB[371] BLB[372] BLB[373]
+ BLB[374] BLB[375] BLB[376] BLB[377] BLB[378] BLB[379] BLB[380] BLB[381]
+ BLB[382] BLB[383] BLB[384] BLB[385] BLB[386] BLB[387] BLB[388] BLB[389]
+ BLB[390] BLB[391] BLB[392] BLB[393] BLB[394] BLB[395] BLB[396] BLB[397]
+ BLB[398] BLB[399] BLB[400] BLB[401] BLB[402] BLB[403] BLB[404] BLB[405]
+ BLB[406] BLB[407] BLB[408] BLB[409] BLB[410] BLB[411] BLB[412] BLB[413]
+ BLB[414] BLB[415] BLB[416] BLB[417] BLB[418] BLB[419] BLB[420] BLB[421]
+ BLB[422] BLB[423] BLB[424] BLB[425] BLB[426] BLB[427] BLB[428] BLB[429]
+ BLB[430] BLB[431] BLB[432] BLB[433] BLB[434] BLB[435] BLB[436] BLB[437]
+ BLB[438] BLB[439] BLB[440] BLB[441] BLB[442] BLB[443] BLB[444] BLB[445]
+ BLB[446] BLB[447] BLB[448] BLB[449] BLB[450] BLB[451] BLB[452] BLB[453]
+ BLB[454] BLB[455] BLB[456] BLB[457] BLB[458] BLB[459] BLB[460] BLB[461]
+ BLB[462] BLB[463] BLB[464] BLB[465] BLB[466] BLB[467] BLB[468] BLB[469]
+ BLB[470] BLB[471] BLB[472] BLB[473] BLB[474] BLB[475] BLB[476] BLB[477]
+ BLB[478] BLB[479] BLB[480] BLB[481] BLB[482] BLB[483] BLB[484] BLB[485]
+ BLB[486] BLB[487] BLB[488] BLB[489] BLB[490] BLB[491] BLB[492] BLB[493]
+ BLB[494] BLB[495] BLB[496] BLB[497] BLB[498] BLB[499] BLB[500] BLB[501]
+ BLB[502] BLB[503] BLB[504] BLB[505] BLB[506] BLB[507] BLB[508] BLB[509]
+ BLB[510] BLB[511] BLB[512] BLB[513] BLB[514] BLB[515] BLB[516] BLB[517]
+ BLB[518] BLB[519] BLB[520] BLB[521] BLB[522] BLB[523] BLB[524] BLB[525]
+ BLB[526] BLB[527] BLB[528] BLB[529] BLB[530] BLB[531] BLB[532] BLB[533]
+ BLB[534] BLB[535] BLB[536] BLB[537] BLB[538] BLB[539] BLB[540] BLB[541]
+ BLB[542] BLB[543] BLB[544] BLB[545] BLB[546] BLB[547] BLB[548] BLB[549]
+ BLB[550] BLB[551] BLB[552] BLB[553] BLB[554] BLB[555] BLB[556] BLB[557]
+ BLB[558] BLB[559] BLB[560] BLB[561] BLB[562] BLB[563] BLB[564] BLB[565]
+ BLB[566] BLB[567] BLB[568] BLB[569] BLB[570] BLB[571] BLB[572] BLB[573]
+ BLB[574] BLB[575] WL[254] WL[255] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22]
+ GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31]
+ GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4]
+ GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13]
+ GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21]
+ GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29]
+ GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_X
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_LIO_L_SD BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3]
+ BLB_DN[4] BLB_DN[5] BLB_DN[6] BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10]
+ BLB_DN[11] BLB_DN[12] BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_DN[16] BLB_DN[17]
+ BLB_DN[18] BLB_DN[19] BLB_DN[20] BLB_DN[21] BLB_DN[22] BLB_DN[23] BLB_DN[24]
+ BLB_DN[25] BLB_DN[26] BLB_DN[27] BLB_DN[28] BLB_DN[29] BLB_DN[30] BLB_DN[31]
+ BLB_DN[32] BLB_DN[33] BLB_DN[34] BLB_DN[35] BLB_DN[36] BLB_DN[37] BLB_DN[38]
+ BLB_DN[39] BLB_DN[40] BLB_DN[41] BLB_DN[42] BLB_DN[43] BLB_DN[44] BLB_DN[45]
+ BLB_DN[46] BLB_DN[47] BLB_DN[48] BLB_DN[49] BLB_DN[50] BLB_DN[51] BLB_DN[52]
+ BLB_DN[53] BLB_DN[54] BLB_DN[55] BLB_DN[56] BLB_DN[57] BLB_DN[58] BLB_DN[59]
+ BLB_DN[60] BLB_DN[61] BLB_DN[62] BLB_DN[63] BLB_DN[64] BLB_DN[65] BLB_DN[66]
+ BLB_DN[67] BLB_DN[68] BLB_DN[69] BLB_DN[70] BLB_DN[71] BLB_DN[72] BLB_DN[73]
+ BLB_DN[74] BLB_DN[75] BLB_DN[76] BLB_DN[77] BLB_DN[78] BLB_DN[79] BLB_DN[80]
+ BLB_DN[81] BLB_DN[82] BLB_DN[83] BLB_DN[84] BLB_DN[85] BLB_DN[86] BLB_DN[87]
+ BLB_DN[88] BLB_DN[89] BLB_DN[90] BLB_DN[91] BLB_DN[92] BLB_DN[93] BLB_DN[94]
+ BLB_DN[95] BLB_DN[96] BLB_DN[97] BLB_DN[98] BLB_DN[99] BLB_DN[100] BLB_DN[101]
+ BLB_DN[102] BLB_DN[103] BLB_DN[104] BLB_DN[105] BLB_DN[106] BLB_DN[107]
+ BLB_DN[108] BLB_DN[109] BLB_DN[110] BLB_DN[111] BLB_DN[112] BLB_DN[113]
+ BLB_DN[114] BLB_DN[115] BLB_DN[116] BLB_DN[117] BLB_DN[118] BLB_DN[119]
+ BLB_DN[120] BLB_DN[121] BLB_DN[122] BLB_DN[123] BLB_DN[124] BLB_DN[125]
+ BLB_DN[126] BLB_DN[127] BLB_DN[128] BLB_DN[129] BLB_DN[130] BLB_DN[131]
+ BLB_DN[132] BLB_DN[133] BLB_DN[134] BLB_DN[135] BLB_DN[136] BLB_DN[137]
+ BLB_DN[138] BLB_DN[139] BLB_DN[140] BLB_DN[141] BLB_DN[142] BLB_DN[143]
+ BLB_DN[144] BLB_DN[145] BLB_DN[146] BLB_DN[147] BLB_DN[148] BLB_DN[149]
+ BLB_DN[150] BLB_DN[151] BLB_DN[152] BLB_DN[153] BLB_DN[154] BLB_DN[155]
+ BLB_DN[156] BLB_DN[157] BLB_DN[158] BLB_DN[159] BLB_DN[160] BLB_DN[161]
+ BLB_DN[162] BLB_DN[163] BLB_DN[164] BLB_DN[165] BLB_DN[166] BLB_DN[167]
+ BLB_DN[168] BLB_DN[169] BLB_DN[170] BLB_DN[171] BLB_DN[172] BLB_DN[173]
+ BLB_DN[174] BLB_DN[175] BLB_DN[176] BLB_DN[177] BLB_DN[178] BLB_DN[179]
+ BLB_DN[180] BLB_DN[181] BLB_DN[182] BLB_DN[183] BLB_DN[184] BLB_DN[185]
+ BLB_DN[186] BLB_DN[187] BLB_DN[188] BLB_DN[189] BLB_DN[190] BLB_DN[191]
+ BLB_DN[192] BLB_DN[193] BLB_DN[194] BLB_DN[195] BLB_DN[196] BLB_DN[197]
+ BLB_DN[198] BLB_DN[199] BLB_DN[200] BLB_DN[201] BLB_DN[202] BLB_DN[203]
+ BLB_DN[204] BLB_DN[205] BLB_DN[206] BLB_DN[207] BLB_DN[208] BLB_DN[209]
+ BLB_DN[210] BLB_DN[211] BLB_DN[212] BLB_DN[213] BLB_DN[214] BLB_DN[215]
+ BLB_DN[216] BLB_DN[217] BLB_DN[218] BLB_DN[219] BLB_DN[220] BLB_DN[221]
+ BLB_DN[222] BLB_DN[223] BLB_DN[224] BLB_DN[225] BLB_DN[226] BLB_DN[227]
+ BLB_DN[228] BLB_DN[229] BLB_DN[230] BLB_DN[231] BLB_DN[232] BLB_DN[233]
+ BLB_DN[234] BLB_DN[235] BLB_DN[236] BLB_DN[237] BLB_DN[238] BLB_DN[239]
+ BLB_DN[240] BLB_DN[241] BLB_DN[242] BLB_DN[243] BLB_DN[244] BLB_DN[245]
+ BLB_DN[246] BLB_DN[247] BLB_DN[248] BLB_DN[249] BLB_DN[250] BLB_DN[251]
+ BLB_DN[252] BLB_DN[253] BLB_DN[254] BLB_DN[255] BLB_DN[256] BLB_DN[257]
+ BLB_DN[258] BLB_DN[259] BLB_DN[260] BLB_DN[261] BLB_DN[262] BLB_DN[263]
+ BLB_DN[264] BLB_DN[265] BLB_DN[266] BLB_DN[267] BLB_DN[268] BLB_DN[269]
+ BLB_DN[270] BLB_DN[271] BLB_DN[272] BLB_DN[273] BLB_DN[274] BLB_DN[275]
+ BLB_DN[276] BLB_DN[277] BLB_DN[278] BLB_DN[279] BLB_DN[280] BLB_DN[281]
+ BLB_DN[282] BLB_DN[283] BLB_DN[284] BLB_DN[285] BLB_DN[286] BLB_DN[287]
+ BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] BLB_UP[4] BLB_UP[5] BLB_UP[6]
+ BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10] BLB_UP[11] BLB_UP[12] BLB_UP[13]
+ BLB_UP[14] BLB_UP[15] BLB_UP[16] BLB_UP[17] BLB_UP[18] BLB_UP[19] BLB_UP[20]
+ BLB_UP[21] BLB_UP[22] BLB_UP[23] BLB_UP[24] BLB_UP[25] BLB_UP[26] BLB_UP[27]
+ BLB_UP[28] BLB_UP[29] BLB_UP[30] BLB_UP[31] BLB_UP[32] BLB_UP[33] BLB_UP[34]
+ BLB_UP[35] BLB_UP[36] BLB_UP[37] BLB_UP[38] BLB_UP[39] BLB_UP[40] BLB_UP[41]
+ BLB_UP[42] BLB_UP[43] BLB_UP[44] BLB_UP[45] BLB_UP[46] BLB_UP[47] BLB_UP[48]
+ BLB_UP[49] BLB_UP[50] BLB_UP[51] BLB_UP[52] BLB_UP[53] BLB_UP[54] BLB_UP[55]
+ BLB_UP[56] BLB_UP[57] BLB_UP[58] BLB_UP[59] BLB_UP[60] BLB_UP[61] BLB_UP[62]
+ BLB_UP[63] BLB_UP[64] BLB_UP[65] BLB_UP[66] BLB_UP[67] BLB_UP[68] BLB_UP[69]
+ BLB_UP[70] BLB_UP[71] BLB_UP[72] BLB_UP[73] BLB_UP[74] BLB_UP[75] BLB_UP[76]
+ BLB_UP[77] BLB_UP[78] BLB_UP[79] BLB_UP[80] BLB_UP[81] BLB_UP[82] BLB_UP[83]
+ BLB_UP[84] BLB_UP[85] BLB_UP[86] BLB_UP[87] BLB_UP[88] BLB_UP[89] BLB_UP[90]
+ BLB_UP[91] BLB_UP[92] BLB_UP[93] BLB_UP[94] BLB_UP[95] BLB_UP[96] BLB_UP[97]
+ BLB_UP[98] BLB_UP[99] BLB_UP[100] BLB_UP[101] BLB_UP[102] BLB_UP[103]
+ BLB_UP[104] BLB_UP[105] BLB_UP[106] BLB_UP[107] BLB_UP[108] BLB_UP[109]
+ BLB_UP[110] BLB_UP[111] BLB_UP[112] BLB_UP[113] BLB_UP[114] BLB_UP[115]
+ BLB_UP[116] BLB_UP[117] BLB_UP[118] BLB_UP[119] BLB_UP[120] BLB_UP[121]
+ BLB_UP[122] BLB_UP[123] BLB_UP[124] BLB_UP[125] BLB_UP[126] BLB_UP[127]
+ BLB_UP[128] BLB_UP[129] BLB_UP[130] BLB_UP[131] BLB_UP[132] BLB_UP[133]
+ BLB_UP[134] BLB_UP[135] BLB_UP[136] BLB_UP[137] BLB_UP[138] BLB_UP[139]
+ BLB_UP[140] BLB_UP[141] BLB_UP[142] BLB_UP[143] BLB_UP[144] BLB_UP[145]
+ BLB_UP[146] BLB_UP[147] BLB_UP[148] BLB_UP[149] BLB_UP[150] BLB_UP[151]
+ BLB_UP[152] BLB_UP[153] BLB_UP[154] BLB_UP[155] BLB_UP[156] BLB_UP[157]
+ BLB_UP[158] BLB_UP[159] BLB_UP[160] BLB_UP[161] BLB_UP[162] BLB_UP[163]
+ BLB_UP[164] BLB_UP[165] BLB_UP[166] BLB_UP[167] BLB_UP[168] BLB_UP[169]
+ BLB_UP[170] BLB_UP[171] BLB_UP[172] BLB_UP[173] BLB_UP[174] BLB_UP[175]
+ BLB_UP[176] BLB_UP[177] BLB_UP[178] BLB_UP[179] BLB_UP[180] BLB_UP[181]
+ BLB_UP[182] BLB_UP[183] BLB_UP[184] BLB_UP[185] BLB_UP[186] BLB_UP[187]
+ BLB_UP[188] BLB_UP[189] BLB_UP[190] BLB_UP[191] BLB_UP[192] BLB_UP[193]
+ BLB_UP[194] BLB_UP[195] BLB_UP[196] BLB_UP[197] BLB_UP[198] BLB_UP[199]
+ BLB_UP[200] BLB_UP[201] BLB_UP[202] BLB_UP[203] BLB_UP[204] BLB_UP[205]
+ BLB_UP[206] BLB_UP[207] BLB_UP[208] BLB_UP[209] BLB_UP[210] BLB_UP[211]
+ BLB_UP[212] BLB_UP[213] BLB_UP[214] BLB_UP[215] BLB_UP[216] BLB_UP[217]
+ BLB_UP[218] BLB_UP[219] BLB_UP[220] BLB_UP[221] BLB_UP[222] BLB_UP[223]
+ BLB_UP[224] BLB_UP[225] BLB_UP[226] BLB_UP[227] BLB_UP[228] BLB_UP[229]
+ BLB_UP[230] BLB_UP[231] BLB_UP[232] BLB_UP[233] BLB_UP[234] BLB_UP[235]
+ BLB_UP[236] BLB_UP[237] BLB_UP[238] BLB_UP[239] BLB_UP[240] BLB_UP[241]
+ BLB_UP[242] BLB_UP[243] BLB_UP[244] BLB_UP[245] BLB_UP[246] BLB_UP[247]
+ BLB_UP[248] BLB_UP[249] BLB_UP[250] BLB_UP[251] BLB_UP[252] BLB_UP[253]
+ BLB_UP[254] BLB_UP[255] BLB_UP[256] BLB_UP[257] BLB_UP[258] BLB_UP[259]
+ BLB_UP[260] BLB_UP[261] BLB_UP[262] BLB_UP[263] BLB_UP[264] BLB_UP[265]
+ BLB_UP[266] BLB_UP[267] BLB_UP[268] BLB_UP[269] BLB_UP[270] BLB_UP[271]
+ BLB_UP[272] BLB_UP[273] BLB_UP[274] BLB_UP[275] BLB_UP[276] BLB_UP[277]
+ BLB_UP[278] BLB_UP[279] BLB_UP[280] BLB_UP[281] BLB_UP[282] BLB_UP[283]
+ BLB_UP[284] BLB_UP[285] BLB_UP[286] BLB_UP[287] BLEQ_DN BLEQ_UP BL_DN[0]
+ BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] BL_DN[8]
+ BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14] BL_DN[15] BL_DN[16]
+ BL_DN[17] BL_DN[18] BL_DN[19] BL_DN[20] BL_DN[21] BL_DN[22] BL_DN[23]
+ BL_DN[24] BL_DN[25] BL_DN[26] BL_DN[27] BL_DN[28] BL_DN[29] BL_DN[30]
+ BL_DN[31] BL_DN[32] BL_DN[33] BL_DN[34] BL_DN[35] BL_DN[36] BL_DN[37]
+ BL_DN[38] BL_DN[39] BL_DN[40] BL_DN[41] BL_DN[42] BL_DN[43] BL_DN[44]
+ BL_DN[45] BL_DN[46] BL_DN[47] BL_DN[48] BL_DN[49] BL_DN[50] BL_DN[51]
+ BL_DN[52] BL_DN[53] BL_DN[54] BL_DN[55] BL_DN[56] BL_DN[57] BL_DN[58]
+ BL_DN[59] BL_DN[60] BL_DN[61] BL_DN[62] BL_DN[63] BL_DN[64] BL_DN[65]
+ BL_DN[66] BL_DN[67] BL_DN[68] BL_DN[69] BL_DN[70] BL_DN[71] BL_DN[72]
+ BL_DN[73] BL_DN[74] BL_DN[75] BL_DN[76] BL_DN[77] BL_DN[78] BL_DN[79]
+ BL_DN[80] BL_DN[81] BL_DN[82] BL_DN[83] BL_DN[84] BL_DN[85] BL_DN[86]
+ BL_DN[87] BL_DN[88] BL_DN[89] BL_DN[90] BL_DN[91] BL_DN[92] BL_DN[93]
+ BL_DN[94] BL_DN[95] BL_DN[96] BL_DN[97] BL_DN[98] BL_DN[99] BL_DN[100]
+ BL_DN[101] BL_DN[102] BL_DN[103] BL_DN[104] BL_DN[105] BL_DN[106] BL_DN[107]
+ BL_DN[108] BL_DN[109] BL_DN[110] BL_DN[111] BL_DN[112] BL_DN[113] BL_DN[114]
+ BL_DN[115] BL_DN[116] BL_DN[117] BL_DN[118] BL_DN[119] BL_DN[120] BL_DN[121]
+ BL_DN[122] BL_DN[123] BL_DN[124] BL_DN[125] BL_DN[126] BL_DN[127] BL_DN[128]
+ BL_DN[129] BL_DN[130] BL_DN[131] BL_DN[132] BL_DN[133] BL_DN[134] BL_DN[135]
+ BL_DN[136] BL_DN[137] BL_DN[138] BL_DN[139] BL_DN[140] BL_DN[141] BL_DN[142]
+ BL_DN[143] BL_DN[144] BL_DN[145] BL_DN[146] BL_DN[147] BL_DN[148] BL_DN[149]
+ BL_DN[150] BL_DN[151] BL_DN[152] BL_DN[153] BL_DN[154] BL_DN[155] BL_DN[156]
+ BL_DN[157] BL_DN[158] BL_DN[159] BL_DN[160] BL_DN[161] BL_DN[162] BL_DN[163]
+ BL_DN[164] BL_DN[165] BL_DN[166] BL_DN[167] BL_DN[168] BL_DN[169] BL_DN[170]
+ BL_DN[171] BL_DN[172] BL_DN[173] BL_DN[174] BL_DN[175] BL_DN[176] BL_DN[177]
+ BL_DN[178] BL_DN[179] BL_DN[180] BL_DN[181] BL_DN[182] BL_DN[183] BL_DN[184]
+ BL_DN[185] BL_DN[186] BL_DN[187] BL_DN[188] BL_DN[189] BL_DN[190] BL_DN[191]
+ BL_DN[192] BL_DN[193] BL_DN[194] BL_DN[195] BL_DN[196] BL_DN[197] BL_DN[198]
+ BL_DN[199] BL_DN[200] BL_DN[201] BL_DN[202] BL_DN[203] BL_DN[204] BL_DN[205]
+ BL_DN[206] BL_DN[207] BL_DN[208] BL_DN[209] BL_DN[210] BL_DN[211] BL_DN[212]
+ BL_DN[213] BL_DN[214] BL_DN[215] BL_DN[216] BL_DN[217] BL_DN[218] BL_DN[219]
+ BL_DN[220] BL_DN[221] BL_DN[222] BL_DN[223] BL_DN[224] BL_DN[225] BL_DN[226]
+ BL_DN[227] BL_DN[228] BL_DN[229] BL_DN[230] BL_DN[231] BL_DN[232] BL_DN[233]
+ BL_DN[234] BL_DN[235] BL_DN[236] BL_DN[237] BL_DN[238] BL_DN[239] BL_DN[240]
+ BL_DN[241] BL_DN[242] BL_DN[243] BL_DN[244] BL_DN[245] BL_DN[246] BL_DN[247]
+ BL_DN[248] BL_DN[249] BL_DN[250] BL_DN[251] BL_DN[252] BL_DN[253] BL_DN[254]
+ BL_DN[255] BL_DN[256] BL_DN[257] BL_DN[258] BL_DN[259] BL_DN[260] BL_DN[261]
+ BL_DN[262] BL_DN[263] BL_DN[264] BL_DN[265] BL_DN[266] BL_DN[267] BL_DN[268]
+ BL_DN[269] BL_DN[270] BL_DN[271] BL_DN[272] BL_DN[273] BL_DN[274] BL_DN[275]
+ BL_DN[276] BL_DN[277] BL_DN[278] BL_DN[279] BL_DN[280] BL_DN[281] BL_DN[282]
+ BL_DN[283] BL_DN[284] BL_DN[285] BL_DN[286] BL_DN[287] BL_UP[0] BL_UP[1]
+ BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] BL_UP[7] BL_UP[8] BL_UP[9]
+ BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14] BL_UP[15] BL_UP[16]
+ BL_UP[17] BL_UP[18] BL_UP[19] BL_UP[20] BL_UP[21] BL_UP[22] BL_UP[23]
+ BL_UP[24] BL_UP[25] BL_UP[26] BL_UP[27] BL_UP[28] BL_UP[29] BL_UP[30]
+ BL_UP[31] BL_UP[32] BL_UP[33] BL_UP[34] BL_UP[35] BL_UP[36] BL_UP[37]
+ BL_UP[38] BL_UP[39] BL_UP[40] BL_UP[41] BL_UP[42] BL_UP[43] BL_UP[44]
+ BL_UP[45] BL_UP[46] BL_UP[47] BL_UP[48] BL_UP[49] BL_UP[50] BL_UP[51]
+ BL_UP[52] BL_UP[53] BL_UP[54] BL_UP[55] BL_UP[56] BL_UP[57] BL_UP[58]
+ BL_UP[59] BL_UP[60] BL_UP[61] BL_UP[62] BL_UP[63] BL_UP[64] BL_UP[65]
+ BL_UP[66] BL_UP[67] BL_UP[68] BL_UP[69] BL_UP[70] BL_UP[71] BL_UP[72]
+ BL_UP[73] BL_UP[74] BL_UP[75] BL_UP[76] BL_UP[77] BL_UP[78] BL_UP[79]
+ BL_UP[80] BL_UP[81] BL_UP[82] BL_UP[83] BL_UP[84] BL_UP[85] BL_UP[86]
+ BL_UP[87] BL_UP[88] BL_UP[89] BL_UP[90] BL_UP[91] BL_UP[92] BL_UP[93]
+ BL_UP[94] BL_UP[95] BL_UP[96] BL_UP[97] BL_UP[98] BL_UP[99] BL_UP[100]
+ BL_UP[101] BL_UP[102] BL_UP[103] BL_UP[104] BL_UP[105] BL_UP[106] BL_UP[107]
+ BL_UP[108] BL_UP[109] BL_UP[110] BL_UP[111] BL_UP[112] BL_UP[113] BL_UP[114]
+ BL_UP[115] BL_UP[116] BL_UP[117] BL_UP[118] BL_UP[119] BL_UP[120] BL_UP[121]
+ BL_UP[122] BL_UP[123] BL_UP[124] BL_UP[125] BL_UP[126] BL_UP[127] BL_UP[128]
+ BL_UP[129] BL_UP[130] BL_UP[131] BL_UP[132] BL_UP[133] BL_UP[134] BL_UP[135]
+ BL_UP[136] BL_UP[137] BL_UP[138] BL_UP[139] BL_UP[140] BL_UP[141] BL_UP[142]
+ BL_UP[143] BL_UP[144] BL_UP[145] BL_UP[146] BL_UP[147] BL_UP[148] BL_UP[149]
+ BL_UP[150] BL_UP[151] BL_UP[152] BL_UP[153] BL_UP[154] BL_UP[155] BL_UP[156]
+ BL_UP[157] BL_UP[158] BL_UP[159] BL_UP[160] BL_UP[161] BL_UP[162] BL_UP[163]
+ BL_UP[164] BL_UP[165] BL_UP[166] BL_UP[167] BL_UP[168] BL_UP[169] BL_UP[170]
+ BL_UP[171] BL_UP[172] BL_UP[173] BL_UP[174] BL_UP[175] BL_UP[176] BL_UP[177]
+ BL_UP[178] BL_UP[179] BL_UP[180] BL_UP[181] BL_UP[182] BL_UP[183] BL_UP[184]
+ BL_UP[185] BL_UP[186] BL_UP[187] BL_UP[188] BL_UP[189] BL_UP[190] BL_UP[191]
+ BL_UP[192] BL_UP[193] BL_UP[194] BL_UP[195] BL_UP[196] BL_UP[197] BL_UP[198]
+ BL_UP[199] BL_UP[200] BL_UP[201] BL_UP[202] BL_UP[203] BL_UP[204] BL_UP[205]
+ BL_UP[206] BL_UP[207] BL_UP[208] BL_UP[209] BL_UP[210] BL_UP[211] BL_UP[212]
+ BL_UP[213] BL_UP[214] BL_UP[215] BL_UP[216] BL_UP[217] BL_UP[218] BL_UP[219]
+ BL_UP[220] BL_UP[221] BL_UP[222] BL_UP[223] BL_UP[224] BL_UP[225] BL_UP[226]
+ BL_UP[227] BL_UP[228] BL_UP[229] BL_UP[230] BL_UP[231] BL_UP[232] BL_UP[233]
+ BL_UP[234] BL_UP[235] BL_UP[236] BL_UP[237] BL_UP[238] BL_UP[239] BL_UP[240]
+ BL_UP[241] BL_UP[242] BL_UP[243] BL_UP[244] BL_UP[245] BL_UP[246] BL_UP[247]
+ BL_UP[248] BL_UP[249] BL_UP[250] BL_UP[251] BL_UP[252] BL_UP[253] BL_UP[254]
+ BL_UP[255] BL_UP[256] BL_UP[257] BL_UP[258] BL_UP[259] BL_UP[260] BL_UP[261]
+ BL_UP[262] BL_UP[263] BL_UP[264] BL_UP[265] BL_UP[266] BL_UP[267] BL_UP[268]
+ BL_UP[269] BL_UP[270] BL_UP[271] BL_UP[272] BL_UP[273] BL_UP[274] BL_UP[275]
+ BL_UP[276] BL_UP[277] BL_UP[278] BL_UP[279] BL_UP[280] BL_UP[281] BL_UP[282]
+ BL_UP[283] BL_UP[284] BL_UP[285] BL_UP[286] BL_UP[287] GBL[0] GBL[1] GBL[2]
+ GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12]
+ GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBLB[0] GBLB[1] GBLB[2] GBLB[3]
+ GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12]
+ GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9]
+ GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] LIOPD PDI PDOX
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
XLIO_M16_SD_0 BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5]
+ BLB_DN[6] BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12]
+ BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3]
+ BLB_UP[4] BLB_UP[5] BLB_UP[6] BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10]
+ BLB_UP[11] BLB_UP[12] BLB_UP[13] BLB_UP[14] BLB_UP[15] BLEQ_DN BLEQ_UP
+ BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7]
+ BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14] BL_DN[15]
+ BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] BL_UP[7]
+ BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14] BL_UP[15]
+ GBL[0] GBLB[0] GW[0] GWB[0] LIOPD PDO1 PDO0 PDO0 RE SAEB VXDDAI VDDI VSSI WE
+ YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6]
+ Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_1 BLB_DN[16] BLB_DN[17] BLB_DN[18] BLB_DN[19] BLB_DN[20] BLB_DN[21]
+ BLB_DN[22] BLB_DN[23] BLB_DN[24] BLB_DN[25] BLB_DN[26] BLB_DN[27] BLB_DN[28]
+ BLB_DN[29] BLB_DN[30] BLB_DN[31] BLB_UP[16] BLB_UP[17] BLB_UP[18] BLB_UP[19]
+ BLB_UP[20] BLB_UP[21] BLB_UP[22] BLB_UP[23] BLB_UP[24] BLB_UP[25] BLB_UP[26]
+ BLB_UP[27] BLB_UP[28] BLB_UP[29] BLB_UP[30] BLB_UP[31] BLEQ_DN BLEQ_UP
+ BL_DN[16] BL_DN[17] BL_DN[18] BL_DN[19] BL_DN[20] BL_DN[21] BL_DN[22]
+ BL_DN[23] BL_DN[24] BL_DN[25] BL_DN[26] BL_DN[27] BL_DN[28] BL_DN[29]
+ BL_DN[30] BL_DN[31] BL_UP[16] BL_UP[17] BL_UP[18] BL_UP[19] BL_UP[20]
+ BL_UP[21] BL_UP[22] BL_UP[23] BL_UP[24] BL_UP[25] BL_UP[26] BL_UP[27]
+ BL_UP[28] BL_UP[29] BL_UP[30] BL_UP[31] GBL[1] GBLB[1] GW[1] GWB[1] LIOPD PDO2
+ PDO1 PDO0 RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1]
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2]
+ Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_2 BLB_DN[32] BLB_DN[33] BLB_DN[34] BLB_DN[35] BLB_DN[36] BLB_DN[37]
+ BLB_DN[38] BLB_DN[39] BLB_DN[40] BLB_DN[41] BLB_DN[42] BLB_DN[43] BLB_DN[44]
+ BLB_DN[45] BLB_DN[46] BLB_DN[47] BLB_UP[32] BLB_UP[33] BLB_UP[34] BLB_UP[35]
+ BLB_UP[36] BLB_UP[37] BLB_UP[38] BLB_UP[39] BLB_UP[40] BLB_UP[41] BLB_UP[42]
+ BLB_UP[43] BLB_UP[44] BLB_UP[45] BLB_UP[46] BLB_UP[47] BLEQ_DN BLEQ_UP
+ BL_DN[32] BL_DN[33] BL_DN[34] BL_DN[35] BL_DN[36] BL_DN[37] BL_DN[38]
+ BL_DN[39] BL_DN[40] BL_DN[41] BL_DN[42] BL_DN[43] BL_DN[44] BL_DN[45]
+ BL_DN[46] BL_DN[47] BL_UP[32] BL_UP[33] BL_UP[34] BL_UP[35] BL_UP[36]
+ BL_UP[37] BL_UP[38] BL_UP[39] BL_UP[40] BL_UP[41] BL_UP[42] BL_UP[43]
+ BL_UP[44] BL_UP[45] BL_UP[46] BL_UP[47] GBL[2] GBLB[2] GW[2] GWB[2] LIOPD PDO3
+ PDO2 PDO0 RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1]
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2]
+ Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_3 BLB_DN[48] BLB_DN[49] BLB_DN[50] BLB_DN[51] BLB_DN[52] BLB_DN[53]
+ BLB_DN[54] BLB_DN[55] BLB_DN[56] BLB_DN[57] BLB_DN[58] BLB_DN[59] BLB_DN[60]
+ BLB_DN[61] BLB_DN[62] BLB_DN[63] BLB_UP[48] BLB_UP[49] BLB_UP[50] BLB_UP[51]
+ BLB_UP[52] BLB_UP[53] BLB_UP[54] BLB_UP[55] BLB_UP[56] BLB_UP[57] BLB_UP[58]
+ BLB_UP[59] BLB_UP[60] BLB_UP[61] BLB_UP[62] BLB_UP[63] BLEQ_DN BLEQ_UP
+ BL_DN[48] BL_DN[49] BL_DN[50] BL_DN[51] BL_DN[52] BL_DN[53] BL_DN[54]
+ BL_DN[55] BL_DN[56] BL_DN[57] BL_DN[58] BL_DN[59] BL_DN[60] BL_DN[61]
+ BL_DN[62] BL_DN[63] BL_UP[48] BL_UP[49] BL_UP[50] BL_UP[51] BL_UP[52]
+ BL_UP[53] BL_UP[54] BL_UP[55] BL_UP[56] BL_UP[57] BL_UP[58] BL_UP[59]
+ BL_UP[60] BL_UP[61] BL_UP[62] BL_UP[63] GBL[3] GBLB[3] GW[3] GWB[3] LIOPD PDO4
+ PDO3 PDO0 RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1]
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2]
+ Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_4 BLB_DN[64] BLB_DN[65] BLB_DN[66] BLB_DN[67] BLB_DN[68] BLB_DN[69]
+ BLB_DN[70] BLB_DN[71] BLB_DN[72] BLB_DN[73] BLB_DN[74] BLB_DN[75] BLB_DN[76]
+ BLB_DN[77] BLB_DN[78] BLB_DN[79] BLB_UP[64] BLB_UP[65] BLB_UP[66] BLB_UP[67]
+ BLB_UP[68] BLB_UP[69] BLB_UP[70] BLB_UP[71] BLB_UP[72] BLB_UP[73] BLB_UP[74]
+ BLB_UP[75] BLB_UP[76] BLB_UP[77] BLB_UP[78] BLB_UP[79] BLEQ_DN BLEQ_UP
+ BL_DN[64] BL_DN[65] BL_DN[66] BL_DN[67] BL_DN[68] BL_DN[69] BL_DN[70]
+ BL_DN[71] BL_DN[72] BL_DN[73] BL_DN[74] BL_DN[75] BL_DN[76] BL_DN[77]
+ BL_DN[78] BL_DN[79] BL_UP[64] BL_UP[65] BL_UP[66] BL_UP[67] BL_UP[68]
+ BL_UP[69] BL_UP[70] BL_UP[71] BL_UP[72] BL_UP[73] BL_UP[74] BL_UP[75]
+ BL_UP[76] BL_UP[77] BL_UP[78] BL_UP[79] GBL[4] GBLB[4] GW[4] GWB[4] LIOPD PDO5
+ PDO4 PDO0 RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1]
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2]
+ Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_5 BLB_DN[80] BLB_DN[81] BLB_DN[82] BLB_DN[83] BLB_DN[84] BLB_DN[85]
+ BLB_DN[86] BLB_DN[87] BLB_DN[88] BLB_DN[89] BLB_DN[90] BLB_DN[91] BLB_DN[92]
+ BLB_DN[93] BLB_DN[94] BLB_DN[95] BLB_UP[80] BLB_UP[81] BLB_UP[82] BLB_UP[83]
+ BLB_UP[84] BLB_UP[85] BLB_UP[86] BLB_UP[87] BLB_UP[88] BLB_UP[89] BLB_UP[90]
+ BLB_UP[91] BLB_UP[92] BLB_UP[93] BLB_UP[94] BLB_UP[95] BLEQ_DN BLEQ_UP
+ BL_DN[80] BL_DN[81] BL_DN[82] BL_DN[83] BL_DN[84] BL_DN[85] BL_DN[86]
+ BL_DN[87] BL_DN[88] BL_DN[89] BL_DN[90] BL_DN[91] BL_DN[92] BL_DN[93]
+ BL_DN[94] BL_DN[95] BL_UP[80] BL_UP[81] BL_UP[82] BL_UP[83] BL_UP[84]
+ BL_UP[85] BL_UP[86] BL_UP[87] BL_UP[88] BL_UP[89] BL_UP[90] BL_UP[91]
+ BL_UP[92] BL_UP[93] BL_UP[94] BL_UP[95] GBL[5] GBLB[5] GW[5] GWB[5] LIOPD PDO6
+ PDO5 PDO0 RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1]
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2]
+ Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_6 BLB_DN[96] BLB_DN[97] BLB_DN[98] BLB_DN[99] BLB_DN[100]
+ BLB_DN[101] BLB_DN[102] BLB_DN[103] BLB_DN[104] BLB_DN[105] BLB_DN[106]
+ BLB_DN[107] BLB_DN[108] BLB_DN[109] BLB_DN[110] BLB_DN[111] BLB_UP[96]
+ BLB_UP[97] BLB_UP[98] BLB_UP[99] BLB_UP[100] BLB_UP[101] BLB_UP[102]
+ BLB_UP[103] BLB_UP[104] BLB_UP[105] BLB_UP[106] BLB_UP[107] BLB_UP[108]
+ BLB_UP[109] BLB_UP[110] BLB_UP[111] BLEQ_DN BLEQ_UP BL_DN[96] BL_DN[97]
+ BL_DN[98] BL_DN[99] BL_DN[100] BL_DN[101] BL_DN[102] BL_DN[103] BL_DN[104]
+ BL_DN[105] BL_DN[106] BL_DN[107] BL_DN[108] BL_DN[109] BL_DN[110] BL_DN[111]
+ BL_UP[96] BL_UP[97] BL_UP[98] BL_UP[99] BL_UP[100] BL_UP[101] BL_UP[102]
+ BL_UP[103] BL_UP[104] BL_UP[105] BL_UP[106] BL_UP[107] BL_UP[108] BL_UP[109]
+ BL_UP[110] BL_UP[111] GBL[6] GBLB[6] GW[6] GWB[6] LIOPD PDO7 PDO6 PDO0 RE SAEB
+ VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_7 BLB_DN[112] BLB_DN[113] BLB_DN[114] BLB_DN[115] BLB_DN[116]
+ BLB_DN[117] BLB_DN[118] BLB_DN[119] BLB_DN[120] BLB_DN[121] BLB_DN[122]
+ BLB_DN[123] BLB_DN[124] BLB_DN[125] BLB_DN[126] BLB_DN[127] BLB_UP[112]
+ BLB_UP[113] BLB_UP[114] BLB_UP[115] BLB_UP[116] BLB_UP[117] BLB_UP[118]
+ BLB_UP[119] BLB_UP[120] BLB_UP[121] BLB_UP[122] BLB_UP[123] BLB_UP[124]
+ BLB_UP[125] BLB_UP[126] BLB_UP[127] BLEQ_DN BLEQ_UP BL_DN[112] BL_DN[113]
+ BL_DN[114] BL_DN[115] BL_DN[116] BL_DN[117] BL_DN[118] BL_DN[119] BL_DN[120]
+ BL_DN[121] BL_DN[122] BL_DN[123] BL_DN[124] BL_DN[125] BL_DN[126] BL_DN[127]
+ BL_UP[112] BL_UP[113] BL_UP[114] BL_UP[115] BL_UP[116] BL_UP[117] BL_UP[118]
+ BL_UP[119] BL_UP[120] BL_UP[121] BL_UP[122] BL_UP[123] BL_UP[124] BL_UP[125]
+ BL_UP[126] BL_UP[127] GBL[7] GBLB[7] GW[7] GWB[7] LIOPD PDO8 PDO7 PDO0 RE SAEB
+ VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_8 BLB_DN[128] BLB_DN[129] BLB_DN[130] BLB_DN[131] BLB_DN[132]
+ BLB_DN[133] BLB_DN[134] BLB_DN[135] BLB_DN[136] BLB_DN[137] BLB_DN[138]
+ BLB_DN[139] BLB_DN[140] BLB_DN[141] BLB_DN[142] BLB_DN[143] BLB_UP[128]
+ BLB_UP[129] BLB_UP[130] BLB_UP[131] BLB_UP[132] BLB_UP[133] BLB_UP[134]
+ BLB_UP[135] BLB_UP[136] BLB_UP[137] BLB_UP[138] BLB_UP[139] BLB_UP[140]
+ BLB_UP[141] BLB_UP[142] BLB_UP[143] BLEQ_DN BLEQ_UP BL_DN[128] BL_DN[129]
+ BL_DN[130] BL_DN[131] BL_DN[132] BL_DN[133] BL_DN[134] BL_DN[135] BL_DN[136]
+ BL_DN[137] BL_DN[138] BL_DN[139] BL_DN[140] BL_DN[141] BL_DN[142] BL_DN[143]
+ BL_UP[128] BL_UP[129] BL_UP[130] BL_UP[131] BL_UP[132] BL_UP[133] BL_UP[134]
+ BL_UP[135] BL_UP[136] BL_UP[137] BL_UP[138] BL_UP[139] BL_UP[140] BL_UP[141]
+ BL_UP[142] BL_UP[143] GBL[8] GBLB[8] GW[8] GWB[8] LIOPD PDO9 PDO8 PDO0 RE SAEB
+ VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_9 BLB_DN[144] BLB_DN[145] BLB_DN[146] BLB_DN[147] BLB_DN[148]
+ BLB_DN[149] BLB_DN[150] BLB_DN[151] BLB_DN[152] BLB_DN[153] BLB_DN[154]
+ BLB_DN[155] BLB_DN[156] BLB_DN[157] BLB_DN[158] BLB_DN[159] BLB_UP[144]
+ BLB_UP[145] BLB_UP[146] BLB_UP[147] BLB_UP[148] BLB_UP[149] BLB_UP[150]
+ BLB_UP[151] BLB_UP[152] BLB_UP[153] BLB_UP[154] BLB_UP[155] BLB_UP[156]
+ BLB_UP[157] BLB_UP[158] BLB_UP[159] BLEQ_DN BLEQ_UP BL_DN[144] BL_DN[145]
+ BL_DN[146] BL_DN[147] BL_DN[148] BL_DN[149] BL_DN[150] BL_DN[151] BL_DN[152]
+ BL_DN[153] BL_DN[154] BL_DN[155] BL_DN[156] BL_DN[157] BL_DN[158] BL_DN[159]
+ BL_UP[144] BL_UP[145] BL_UP[146] BL_UP[147] BL_UP[148] BL_UP[149] BL_UP[150]
+ BL_UP[151] BL_UP[152] BL_UP[153] BL_UP[154] BL_UP[155] BL_UP[156] BL_UP[157]
+ BL_UP[158] BL_UP[159] GBL[9] GBLB[9] GW[9] GWB[9] LIOPD PDO10 PDO9 PDO0 RE
+ SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_10 BLB_DN[160] BLB_DN[161] BLB_DN[162] BLB_DN[163] BLB_DN[164]
+ BLB_DN[165] BLB_DN[166] BLB_DN[167] BLB_DN[168] BLB_DN[169] BLB_DN[170]
+ BLB_DN[171] BLB_DN[172] BLB_DN[173] BLB_DN[174] BLB_DN[175] BLB_UP[160]
+ BLB_UP[161] BLB_UP[162] BLB_UP[163] BLB_UP[164] BLB_UP[165] BLB_UP[166]
+ BLB_UP[167] BLB_UP[168] BLB_UP[169] BLB_UP[170] BLB_UP[171] BLB_UP[172]
+ BLB_UP[173] BLB_UP[174] BLB_UP[175] BLEQ_DN BLEQ_UP BL_DN[160] BL_DN[161]
+ BL_DN[162] BL_DN[163] BL_DN[164] BL_DN[165] BL_DN[166] BL_DN[167] BL_DN[168]
+ BL_DN[169] BL_DN[170] BL_DN[171] BL_DN[172] BL_DN[173] BL_DN[174] BL_DN[175]
+ BL_UP[160] BL_UP[161] BL_UP[162] BL_UP[163] BL_UP[164] BL_UP[165] BL_UP[166]
+ BL_UP[167] BL_UP[168] BL_UP[169] BL_UP[170] BL_UP[171] BL_UP[172] BL_UP[173]
+ BL_UP[174] BL_UP[175] GBL[10] GBLB[10] GW[10] GWB[10] LIOPD PDO11 PDO10 PDO0
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_11 BLB_DN[176] BLB_DN[177] BLB_DN[178] BLB_DN[179] BLB_DN[180]
+ BLB_DN[181] BLB_DN[182] BLB_DN[183] BLB_DN[184] BLB_DN[185] BLB_DN[186]
+ BLB_DN[187] BLB_DN[188] BLB_DN[189] BLB_DN[190] BLB_DN[191] BLB_UP[176]
+ BLB_UP[177] BLB_UP[178] BLB_UP[179] BLB_UP[180] BLB_UP[181] BLB_UP[182]
+ BLB_UP[183] BLB_UP[184] BLB_UP[185] BLB_UP[186] BLB_UP[187] BLB_UP[188]
+ BLB_UP[189] BLB_UP[190] BLB_UP[191] BLEQ_DN BLEQ_UP BL_DN[176] BL_DN[177]
+ BL_DN[178] BL_DN[179] BL_DN[180] BL_DN[181] BL_DN[182] BL_DN[183] BL_DN[184]
+ BL_DN[185] BL_DN[186] BL_DN[187] BL_DN[188] BL_DN[189] BL_DN[190] BL_DN[191]
+ BL_UP[176] BL_UP[177] BL_UP[178] BL_UP[179] BL_UP[180] BL_UP[181] BL_UP[182]
+ BL_UP[183] BL_UP[184] BL_UP[185] BL_UP[186] BL_UP[187] BL_UP[188] BL_UP[189]
+ BL_UP[190] BL_UP[191] GBL[11] GBLB[11] GW[11] GWB[11] LIOPD PDO12 PDO11 PDO0
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_12 BLB_DN[192] BLB_DN[193] BLB_DN[194] BLB_DN[195] BLB_DN[196]
+ BLB_DN[197] BLB_DN[198] BLB_DN[199] BLB_DN[200] BLB_DN[201] BLB_DN[202]
+ BLB_DN[203] BLB_DN[204] BLB_DN[205] BLB_DN[206] BLB_DN[207] BLB_UP[192]
+ BLB_UP[193] BLB_UP[194] BLB_UP[195] BLB_UP[196] BLB_UP[197] BLB_UP[198]
+ BLB_UP[199] BLB_UP[200] BLB_UP[201] BLB_UP[202] BLB_UP[203] BLB_UP[204]
+ BLB_UP[205] BLB_UP[206] BLB_UP[207] BLEQ_DN BLEQ_UP BL_DN[192] BL_DN[193]
+ BL_DN[194] BL_DN[195] BL_DN[196] BL_DN[197] BL_DN[198] BL_DN[199] BL_DN[200]
+ BL_DN[201] BL_DN[202] BL_DN[203] BL_DN[204] BL_DN[205] BL_DN[206] BL_DN[207]
+ BL_UP[192] BL_UP[193] BL_UP[194] BL_UP[195] BL_UP[196] BL_UP[197] BL_UP[198]
+ BL_UP[199] BL_UP[200] BL_UP[201] BL_UP[202] BL_UP[203] BL_UP[204] BL_UP[205]
+ BL_UP[206] BL_UP[207] GBL[12] GBLB[12] GW[12] GWB[12] LIOPD PDO13 PDO12 PDO0
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_13 BLB_DN[208] BLB_DN[209] BLB_DN[210] BLB_DN[211] BLB_DN[212]
+ BLB_DN[213] BLB_DN[214] BLB_DN[215] BLB_DN[216] BLB_DN[217] BLB_DN[218]
+ BLB_DN[219] BLB_DN[220] BLB_DN[221] BLB_DN[222] BLB_DN[223] BLB_UP[208]
+ BLB_UP[209] BLB_UP[210] BLB_UP[211] BLB_UP[212] BLB_UP[213] BLB_UP[214]
+ BLB_UP[215] BLB_UP[216] BLB_UP[217] BLB_UP[218] BLB_UP[219] BLB_UP[220]
+ BLB_UP[221] BLB_UP[222] BLB_UP[223] BLEQ_DN BLEQ_UP BL_DN[208] BL_DN[209]
+ BL_DN[210] BL_DN[211] BL_DN[212] BL_DN[213] BL_DN[214] BL_DN[215] BL_DN[216]
+ BL_DN[217] BL_DN[218] BL_DN[219] BL_DN[220] BL_DN[221] BL_DN[222] BL_DN[223]
+ BL_UP[208] BL_UP[209] BL_UP[210] BL_UP[211] BL_UP[212] BL_UP[213] BL_UP[214]
+ BL_UP[215] BL_UP[216] BL_UP[217] BL_UP[218] BL_UP[219] BL_UP[220] BL_UP[221]
+ BL_UP[222] BL_UP[223] GBL[13] GBLB[13] GW[13] GWB[13] LIOPD PDO14 PDO13 PDO0
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_14 BLB_DN[224] BLB_DN[225] BLB_DN[226] BLB_DN[227] BLB_DN[228]
+ BLB_DN[229] BLB_DN[230] BLB_DN[231] BLB_DN[232] BLB_DN[233] BLB_DN[234]
+ BLB_DN[235] BLB_DN[236] BLB_DN[237] BLB_DN[238] BLB_DN[239] BLB_UP[224]
+ BLB_UP[225] BLB_UP[226] BLB_UP[227] BLB_UP[228] BLB_UP[229] BLB_UP[230]
+ BLB_UP[231] BLB_UP[232] BLB_UP[233] BLB_UP[234] BLB_UP[235] BLB_UP[236]
+ BLB_UP[237] BLB_UP[238] BLB_UP[239] BLEQ_DN BLEQ_UP BL_DN[224] BL_DN[225]
+ BL_DN[226] BL_DN[227] BL_DN[228] BL_DN[229] BL_DN[230] BL_DN[231] BL_DN[232]
+ BL_DN[233] BL_DN[234] BL_DN[235] BL_DN[236] BL_DN[237] BL_DN[238] BL_DN[239]
+ BL_UP[224] BL_UP[225] BL_UP[226] BL_UP[227] BL_UP[228] BL_UP[229] BL_UP[230]
+ BL_UP[231] BL_UP[232] BL_UP[233] BL_UP[234] BL_UP[235] BL_UP[236] BL_UP[237]
+ BL_UP[238] BL_UP[239] GBL[14] GBLB[14] GW[14] GWB[14] LIOPD PDO15 PDO14 PDO0
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_15 BLB_DN[240] BLB_DN[241] BLB_DN[242] BLB_DN[243] BLB_DN[244]
+ BLB_DN[245] BLB_DN[246] BLB_DN[247] BLB_DN[248] BLB_DN[249] BLB_DN[250]
+ BLB_DN[251] BLB_DN[252] BLB_DN[253] BLB_DN[254] BLB_DN[255] BLB_UP[240]
+ BLB_UP[241] BLB_UP[242] BLB_UP[243] BLB_UP[244] BLB_UP[245] BLB_UP[246]
+ BLB_UP[247] BLB_UP[248] BLB_UP[249] BLB_UP[250] BLB_UP[251] BLB_UP[252]
+ BLB_UP[253] BLB_UP[254] BLB_UP[255] BLEQ_DN BLEQ_UP BL_DN[240] BL_DN[241]
+ BL_DN[242] BL_DN[243] BL_DN[244] BL_DN[245] BL_DN[246] BL_DN[247] BL_DN[248]
+ BL_DN[249] BL_DN[250] BL_DN[251] BL_DN[252] BL_DN[253] BL_DN[254] BL_DN[255]
+ BL_UP[240] BL_UP[241] BL_UP[242] BL_UP[243] BL_UP[244] BL_UP[245] BL_UP[246]
+ BL_UP[247] BL_UP[248] BL_UP[249] BL_UP[250] BL_UP[251] BL_UP[252] BL_UP[253]
+ BL_UP[254] BL_UP[255] GBL[15] GBLB[15] GW[15] GWB[15] LIOPD PDO16 PDO15 PDO0
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_16 BLB_DN[256] BLB_DN[257] BLB_DN[258] BLB_DN[259] BLB_DN[260]
+ BLB_DN[261] BLB_DN[262] BLB_DN[263] BLB_DN[264] BLB_DN[265] BLB_DN[266]
+ BLB_DN[267] BLB_DN[268] BLB_DN[269] BLB_DN[270] BLB_DN[271] BLB_UP[256]
+ BLB_UP[257] BLB_UP[258] BLB_UP[259] BLB_UP[260] BLB_UP[261] BLB_UP[262]
+ BLB_UP[263] BLB_UP[264] BLB_UP[265] BLB_UP[266] BLB_UP[267] BLB_UP[268]
+ BLB_UP[269] BLB_UP[270] BLB_UP[271] BLEQ_DN BLEQ_UP BL_DN[256] BL_DN[257]
+ BL_DN[258] BL_DN[259] BL_DN[260] BL_DN[261] BL_DN[262] BL_DN[263] BL_DN[264]
+ BL_DN[265] BL_DN[266] BL_DN[267] BL_DN[268] BL_DN[269] BL_DN[270] BL_DN[271]
+ BL_UP[256] BL_UP[257] BL_UP[258] BL_UP[259] BL_UP[260] BL_UP[261] BL_UP[262]
+ BL_UP[263] BL_UP[264] BL_UP[265] BL_UP[266] BL_UP[267] BL_UP[268] BL_UP[269]
+ BL_UP[270] BL_UP[271] GBL[16] GBLB[16] GW[16] GWB[16] LIOPD PDO17 PDO16 PDO0
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_17 BLB_DN[272] BLB_DN[273] BLB_DN[274] BLB_DN[275] BLB_DN[276]
+ BLB_DN[277] BLB_DN[278] BLB_DN[279] BLB_DN[280] BLB_DN[281] BLB_DN[282]
+ BLB_DN[283] BLB_DN[284] BLB_DN[285] BLB_DN[286] BLB_DN[287] BLB_UP[272]
+ BLB_UP[273] BLB_UP[274] BLB_UP[275] BLB_UP[276] BLB_UP[277] BLB_UP[278]
+ BLB_UP[279] BLB_UP[280] BLB_UP[281] BLB_UP[282] BLB_UP[283] BLB_UP[284]
+ BLB_UP[285] BLB_UP[286] BLB_UP[287] BLEQ_DN BLEQ_UP BL_DN[272] BL_DN[273]
+ BL_DN[274] BL_DN[275] BL_DN[276] BL_DN[277] BL_DN[278] BL_DN[279] BL_DN[280]
+ BL_DN[281] BL_DN[282] BL_DN[283] BL_DN[284] BL_DN[285] BL_DN[286] BL_DN[287]
+ BL_UP[272] BL_UP[273] BL_UP[274] BL_UP[275] BL_UP[276] BL_UP[277] BL_UP[278]
+ BL_UP[279] BL_UP[280] BL_UP[281] BL_UP[282] BL_UP[283] BL_UP[284] BL_UP[285]
+ BL_UP[286] BL_UP[287] GBL[17] GBLB[17] GW[17] GWB[17] LIOPD LIOPD PDO17 PDO0
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_LIO_R_SD BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3]
+ BLB_DN[4] BLB_DN[5] BLB_DN[6] BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10]
+ BLB_DN[11] BLB_DN[12] BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_DN[16] BLB_DN[17]
+ BLB_DN[18] BLB_DN[19] BLB_DN[20] BLB_DN[21] BLB_DN[22] BLB_DN[23] BLB_DN[24]
+ BLB_DN[25] BLB_DN[26] BLB_DN[27] BLB_DN[28] BLB_DN[29] BLB_DN[30] BLB_DN[31]
+ BLB_DN[32] BLB_DN[33] BLB_DN[34] BLB_DN[35] BLB_DN[36] BLB_DN[37] BLB_DN[38]
+ BLB_DN[39] BLB_DN[40] BLB_DN[41] BLB_DN[42] BLB_DN[43] BLB_DN[44] BLB_DN[45]
+ BLB_DN[46] BLB_DN[47] BLB_DN[48] BLB_DN[49] BLB_DN[50] BLB_DN[51] BLB_DN[52]
+ BLB_DN[53] BLB_DN[54] BLB_DN[55] BLB_DN[56] BLB_DN[57] BLB_DN[58] BLB_DN[59]
+ BLB_DN[60] BLB_DN[61] BLB_DN[62] BLB_DN[63] BLB_DN[64] BLB_DN[65] BLB_DN[66]
+ BLB_DN[67] BLB_DN[68] BLB_DN[69] BLB_DN[70] BLB_DN[71] BLB_DN[72] BLB_DN[73]
+ BLB_DN[74] BLB_DN[75] BLB_DN[76] BLB_DN[77] BLB_DN[78] BLB_DN[79] BLB_DN[80]
+ BLB_DN[81] BLB_DN[82] BLB_DN[83] BLB_DN[84] BLB_DN[85] BLB_DN[86] BLB_DN[87]
+ BLB_DN[88] BLB_DN[89] BLB_DN[90] BLB_DN[91] BLB_DN[92] BLB_DN[93] BLB_DN[94]
+ BLB_DN[95] BLB_DN[96] BLB_DN[97] BLB_DN[98] BLB_DN[99] BLB_DN[100] BLB_DN[101]
+ BLB_DN[102] BLB_DN[103] BLB_DN[104] BLB_DN[105] BLB_DN[106] BLB_DN[107]
+ BLB_DN[108] BLB_DN[109] BLB_DN[110] BLB_DN[111] BLB_DN[112] BLB_DN[113]
+ BLB_DN[114] BLB_DN[115] BLB_DN[116] BLB_DN[117] BLB_DN[118] BLB_DN[119]
+ BLB_DN[120] BLB_DN[121] BLB_DN[122] BLB_DN[123] BLB_DN[124] BLB_DN[125]
+ BLB_DN[126] BLB_DN[127] BLB_DN[128] BLB_DN[129] BLB_DN[130] BLB_DN[131]
+ BLB_DN[132] BLB_DN[133] BLB_DN[134] BLB_DN[135] BLB_DN[136] BLB_DN[137]
+ BLB_DN[138] BLB_DN[139] BLB_DN[140] BLB_DN[141] BLB_DN[142] BLB_DN[143]
+ BLB_DN[144] BLB_DN[145] BLB_DN[146] BLB_DN[147] BLB_DN[148] BLB_DN[149]
+ BLB_DN[150] BLB_DN[151] BLB_DN[152] BLB_DN[153] BLB_DN[154] BLB_DN[155]
+ BLB_DN[156] BLB_DN[157] BLB_DN[158] BLB_DN[159] BLB_DN[160] BLB_DN[161]
+ BLB_DN[162] BLB_DN[163] BLB_DN[164] BLB_DN[165] BLB_DN[166] BLB_DN[167]
+ BLB_DN[168] BLB_DN[169] BLB_DN[170] BLB_DN[171] BLB_DN[172] BLB_DN[173]
+ BLB_DN[174] BLB_DN[175] BLB_DN[176] BLB_DN[177] BLB_DN[178] BLB_DN[179]
+ BLB_DN[180] BLB_DN[181] BLB_DN[182] BLB_DN[183] BLB_DN[184] BLB_DN[185]
+ BLB_DN[186] BLB_DN[187] BLB_DN[188] BLB_DN[189] BLB_DN[190] BLB_DN[191]
+ BLB_DN[192] BLB_DN[193] BLB_DN[194] BLB_DN[195] BLB_DN[196] BLB_DN[197]
+ BLB_DN[198] BLB_DN[199] BLB_DN[200] BLB_DN[201] BLB_DN[202] BLB_DN[203]
+ BLB_DN[204] BLB_DN[205] BLB_DN[206] BLB_DN[207] BLB_DN[208] BLB_DN[209]
+ BLB_DN[210] BLB_DN[211] BLB_DN[212] BLB_DN[213] BLB_DN[214] BLB_DN[215]
+ BLB_DN[216] BLB_DN[217] BLB_DN[218] BLB_DN[219] BLB_DN[220] BLB_DN[221]
+ BLB_DN[222] BLB_DN[223] BLB_DN[224] BLB_DN[225] BLB_DN[226] BLB_DN[227]
+ BLB_DN[228] BLB_DN[229] BLB_DN[230] BLB_DN[231] BLB_DN[232] BLB_DN[233]
+ BLB_DN[234] BLB_DN[235] BLB_DN[236] BLB_DN[237] BLB_DN[238] BLB_DN[239]
+ BLB_DN[240] BLB_DN[241] BLB_DN[242] BLB_DN[243] BLB_DN[244] BLB_DN[245]
+ BLB_DN[246] BLB_DN[247] BLB_DN[248] BLB_DN[249] BLB_DN[250] BLB_DN[251]
+ BLB_DN[252] BLB_DN[253] BLB_DN[254] BLB_DN[255] BLB_DN[256] BLB_DN[257]
+ BLB_DN[258] BLB_DN[259] BLB_DN[260] BLB_DN[261] BLB_DN[262] BLB_DN[263]
+ BLB_DN[264] BLB_DN[265] BLB_DN[266] BLB_DN[267] BLB_DN[268] BLB_DN[269]
+ BLB_DN[270] BLB_DN[271] BLB_DN[272] BLB_DN[273] BLB_DN[274] BLB_DN[275]
+ BLB_DN[276] BLB_DN[277] BLB_DN[278] BLB_DN[279] BLB_DN[280] BLB_DN[281]
+ BLB_DN[282] BLB_DN[283] BLB_DN[284] BLB_DN[285] BLB_DN[286] BLB_DN[287]
+ BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] BLB_UP[4] BLB_UP[5] BLB_UP[6]
+ BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10] BLB_UP[11] BLB_UP[12] BLB_UP[13]
+ BLB_UP[14] BLB_UP[15] BLB_UP[16] BLB_UP[17] BLB_UP[18] BLB_UP[19] BLB_UP[20]
+ BLB_UP[21] BLB_UP[22] BLB_UP[23] BLB_UP[24] BLB_UP[25] BLB_UP[26] BLB_UP[27]
+ BLB_UP[28] BLB_UP[29] BLB_UP[30] BLB_UP[31] BLB_UP[32] BLB_UP[33] BLB_UP[34]
+ BLB_UP[35] BLB_UP[36] BLB_UP[37] BLB_UP[38] BLB_UP[39] BLB_UP[40] BLB_UP[41]
+ BLB_UP[42] BLB_UP[43] BLB_UP[44] BLB_UP[45] BLB_UP[46] BLB_UP[47] BLB_UP[48]
+ BLB_UP[49] BLB_UP[50] BLB_UP[51] BLB_UP[52] BLB_UP[53] BLB_UP[54] BLB_UP[55]
+ BLB_UP[56] BLB_UP[57] BLB_UP[58] BLB_UP[59] BLB_UP[60] BLB_UP[61] BLB_UP[62]
+ BLB_UP[63] BLB_UP[64] BLB_UP[65] BLB_UP[66] BLB_UP[67] BLB_UP[68] BLB_UP[69]
+ BLB_UP[70] BLB_UP[71] BLB_UP[72] BLB_UP[73] BLB_UP[74] BLB_UP[75] BLB_UP[76]
+ BLB_UP[77] BLB_UP[78] BLB_UP[79] BLB_UP[80] BLB_UP[81] BLB_UP[82] BLB_UP[83]
+ BLB_UP[84] BLB_UP[85] BLB_UP[86] BLB_UP[87] BLB_UP[88] BLB_UP[89] BLB_UP[90]
+ BLB_UP[91] BLB_UP[92] BLB_UP[93] BLB_UP[94] BLB_UP[95] BLB_UP[96] BLB_UP[97]
+ BLB_UP[98] BLB_UP[99] BLB_UP[100] BLB_UP[101] BLB_UP[102] BLB_UP[103]
+ BLB_UP[104] BLB_UP[105] BLB_UP[106] BLB_UP[107] BLB_UP[108] BLB_UP[109]
+ BLB_UP[110] BLB_UP[111] BLB_UP[112] BLB_UP[113] BLB_UP[114] BLB_UP[115]
+ BLB_UP[116] BLB_UP[117] BLB_UP[118] BLB_UP[119] BLB_UP[120] BLB_UP[121]
+ BLB_UP[122] BLB_UP[123] BLB_UP[124] BLB_UP[125] BLB_UP[126] BLB_UP[127]
+ BLB_UP[128] BLB_UP[129] BLB_UP[130] BLB_UP[131] BLB_UP[132] BLB_UP[133]
+ BLB_UP[134] BLB_UP[135] BLB_UP[136] BLB_UP[137] BLB_UP[138] BLB_UP[139]
+ BLB_UP[140] BLB_UP[141] BLB_UP[142] BLB_UP[143] BLB_UP[144] BLB_UP[145]
+ BLB_UP[146] BLB_UP[147] BLB_UP[148] BLB_UP[149] BLB_UP[150] BLB_UP[151]
+ BLB_UP[152] BLB_UP[153] BLB_UP[154] BLB_UP[155] BLB_UP[156] BLB_UP[157]
+ BLB_UP[158] BLB_UP[159] BLB_UP[160] BLB_UP[161] BLB_UP[162] BLB_UP[163]
+ BLB_UP[164] BLB_UP[165] BLB_UP[166] BLB_UP[167] BLB_UP[168] BLB_UP[169]
+ BLB_UP[170] BLB_UP[171] BLB_UP[172] BLB_UP[173] BLB_UP[174] BLB_UP[175]
+ BLB_UP[176] BLB_UP[177] BLB_UP[178] BLB_UP[179] BLB_UP[180] BLB_UP[181]
+ BLB_UP[182] BLB_UP[183] BLB_UP[184] BLB_UP[185] BLB_UP[186] BLB_UP[187]
+ BLB_UP[188] BLB_UP[189] BLB_UP[190] BLB_UP[191] BLB_UP[192] BLB_UP[193]
+ BLB_UP[194] BLB_UP[195] BLB_UP[196] BLB_UP[197] BLB_UP[198] BLB_UP[199]
+ BLB_UP[200] BLB_UP[201] BLB_UP[202] BLB_UP[203] BLB_UP[204] BLB_UP[205]
+ BLB_UP[206] BLB_UP[207] BLB_UP[208] BLB_UP[209] BLB_UP[210] BLB_UP[211]
+ BLB_UP[212] BLB_UP[213] BLB_UP[214] BLB_UP[215] BLB_UP[216] BLB_UP[217]
+ BLB_UP[218] BLB_UP[219] BLB_UP[220] BLB_UP[221] BLB_UP[222] BLB_UP[223]
+ BLB_UP[224] BLB_UP[225] BLB_UP[226] BLB_UP[227] BLB_UP[228] BLB_UP[229]
+ BLB_UP[230] BLB_UP[231] BLB_UP[232] BLB_UP[233] BLB_UP[234] BLB_UP[235]
+ BLB_UP[236] BLB_UP[237] BLB_UP[238] BLB_UP[239] BLB_UP[240] BLB_UP[241]
+ BLB_UP[242] BLB_UP[243] BLB_UP[244] BLB_UP[245] BLB_UP[246] BLB_UP[247]
+ BLB_UP[248] BLB_UP[249] BLB_UP[250] BLB_UP[251] BLB_UP[252] BLB_UP[253]
+ BLB_UP[254] BLB_UP[255] BLB_UP[256] BLB_UP[257] BLB_UP[258] BLB_UP[259]
+ BLB_UP[260] BLB_UP[261] BLB_UP[262] BLB_UP[263] BLB_UP[264] BLB_UP[265]
+ BLB_UP[266] BLB_UP[267] BLB_UP[268] BLB_UP[269] BLB_UP[270] BLB_UP[271]
+ BLB_UP[272] BLB_UP[273] BLB_UP[274] BLB_UP[275] BLB_UP[276] BLB_UP[277]
+ BLB_UP[278] BLB_UP[279] BLB_UP[280] BLB_UP[281] BLB_UP[282] BLB_UP[283]
+ BLB_UP[284] BLB_UP[285] BLB_UP[286] BLB_UP[287] BLEQ_DN BLEQ_UP BL_DN[0]
+ BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] BL_DN[8]
+ BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14] BL_DN[15] BL_DN[16]
+ BL_DN[17] BL_DN[18] BL_DN[19] BL_DN[20] BL_DN[21] BL_DN[22] BL_DN[23]
+ BL_DN[24] BL_DN[25] BL_DN[26] BL_DN[27] BL_DN[28] BL_DN[29] BL_DN[30]
+ BL_DN[31] BL_DN[32] BL_DN[33] BL_DN[34] BL_DN[35] BL_DN[36] BL_DN[37]
+ BL_DN[38] BL_DN[39] BL_DN[40] BL_DN[41] BL_DN[42] BL_DN[43] BL_DN[44]
+ BL_DN[45] BL_DN[46] BL_DN[47] BL_DN[48] BL_DN[49] BL_DN[50] BL_DN[51]
+ BL_DN[52] BL_DN[53] BL_DN[54] BL_DN[55] BL_DN[56] BL_DN[57] BL_DN[58]
+ BL_DN[59] BL_DN[60] BL_DN[61] BL_DN[62] BL_DN[63] BL_DN[64] BL_DN[65]
+ BL_DN[66] BL_DN[67] BL_DN[68] BL_DN[69] BL_DN[70] BL_DN[71] BL_DN[72]
+ BL_DN[73] BL_DN[74] BL_DN[75] BL_DN[76] BL_DN[77] BL_DN[78] BL_DN[79]
+ BL_DN[80] BL_DN[81] BL_DN[82] BL_DN[83] BL_DN[84] BL_DN[85] BL_DN[86]
+ BL_DN[87] BL_DN[88] BL_DN[89] BL_DN[90] BL_DN[91] BL_DN[92] BL_DN[93]
+ BL_DN[94] BL_DN[95] BL_DN[96] BL_DN[97] BL_DN[98] BL_DN[99] BL_DN[100]
+ BL_DN[101] BL_DN[102] BL_DN[103] BL_DN[104] BL_DN[105] BL_DN[106] BL_DN[107]
+ BL_DN[108] BL_DN[109] BL_DN[110] BL_DN[111] BL_DN[112] BL_DN[113] BL_DN[114]
+ BL_DN[115] BL_DN[116] BL_DN[117] BL_DN[118] BL_DN[119] BL_DN[120] BL_DN[121]
+ BL_DN[122] BL_DN[123] BL_DN[124] BL_DN[125] BL_DN[126] BL_DN[127] BL_DN[128]
+ BL_DN[129] BL_DN[130] BL_DN[131] BL_DN[132] BL_DN[133] BL_DN[134] BL_DN[135]
+ BL_DN[136] BL_DN[137] BL_DN[138] BL_DN[139] BL_DN[140] BL_DN[141] BL_DN[142]
+ BL_DN[143] BL_DN[144] BL_DN[145] BL_DN[146] BL_DN[147] BL_DN[148] BL_DN[149]
+ BL_DN[150] BL_DN[151] BL_DN[152] BL_DN[153] BL_DN[154] BL_DN[155] BL_DN[156]
+ BL_DN[157] BL_DN[158] BL_DN[159] BL_DN[160] BL_DN[161] BL_DN[162] BL_DN[163]
+ BL_DN[164] BL_DN[165] BL_DN[166] BL_DN[167] BL_DN[168] BL_DN[169] BL_DN[170]
+ BL_DN[171] BL_DN[172] BL_DN[173] BL_DN[174] BL_DN[175] BL_DN[176] BL_DN[177]
+ BL_DN[178] BL_DN[179] BL_DN[180] BL_DN[181] BL_DN[182] BL_DN[183] BL_DN[184]
+ BL_DN[185] BL_DN[186] BL_DN[187] BL_DN[188] BL_DN[189] BL_DN[190] BL_DN[191]
+ BL_DN[192] BL_DN[193] BL_DN[194] BL_DN[195] BL_DN[196] BL_DN[197] BL_DN[198]
+ BL_DN[199] BL_DN[200] BL_DN[201] BL_DN[202] BL_DN[203] BL_DN[204] BL_DN[205]
+ BL_DN[206] BL_DN[207] BL_DN[208] BL_DN[209] BL_DN[210] BL_DN[211] BL_DN[212]
+ BL_DN[213] BL_DN[214] BL_DN[215] BL_DN[216] BL_DN[217] BL_DN[218] BL_DN[219]
+ BL_DN[220] BL_DN[221] BL_DN[222] BL_DN[223] BL_DN[224] BL_DN[225] BL_DN[226]
+ BL_DN[227] BL_DN[228] BL_DN[229] BL_DN[230] BL_DN[231] BL_DN[232] BL_DN[233]
+ BL_DN[234] BL_DN[235] BL_DN[236] BL_DN[237] BL_DN[238] BL_DN[239] BL_DN[240]
+ BL_DN[241] BL_DN[242] BL_DN[243] BL_DN[244] BL_DN[245] BL_DN[246] BL_DN[247]
+ BL_DN[248] BL_DN[249] BL_DN[250] BL_DN[251] BL_DN[252] BL_DN[253] BL_DN[254]
+ BL_DN[255] BL_DN[256] BL_DN[257] BL_DN[258] BL_DN[259] BL_DN[260] BL_DN[261]
+ BL_DN[262] BL_DN[263] BL_DN[264] BL_DN[265] BL_DN[266] BL_DN[267] BL_DN[268]
+ BL_DN[269] BL_DN[270] BL_DN[271] BL_DN[272] BL_DN[273] BL_DN[274] BL_DN[275]
+ BL_DN[276] BL_DN[277] BL_DN[278] BL_DN[279] BL_DN[280] BL_DN[281] BL_DN[282]
+ BL_DN[283] BL_DN[284] BL_DN[285] BL_DN[286] BL_DN[287] BL_UP[0] BL_UP[1]
+ BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] BL_UP[7] BL_UP[8] BL_UP[9]
+ BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14] BL_UP[15] BL_UP[16]
+ BL_UP[17] BL_UP[18] BL_UP[19] BL_UP[20] BL_UP[21] BL_UP[22] BL_UP[23]
+ BL_UP[24] BL_UP[25] BL_UP[26] BL_UP[27] BL_UP[28] BL_UP[29] BL_UP[30]
+ BL_UP[31] BL_UP[32] BL_UP[33] BL_UP[34] BL_UP[35] BL_UP[36] BL_UP[37]
+ BL_UP[38] BL_UP[39] BL_UP[40] BL_UP[41] BL_UP[42] BL_UP[43] BL_UP[44]
+ BL_UP[45] BL_UP[46] BL_UP[47] BL_UP[48] BL_UP[49] BL_UP[50] BL_UP[51]
+ BL_UP[52] BL_UP[53] BL_UP[54] BL_UP[55] BL_UP[56] BL_UP[57] BL_UP[58]
+ BL_UP[59] BL_UP[60] BL_UP[61] BL_UP[62] BL_UP[63] BL_UP[64] BL_UP[65]
+ BL_UP[66] BL_UP[67] BL_UP[68] BL_UP[69] BL_UP[70] BL_UP[71] BL_UP[72]
+ BL_UP[73] BL_UP[74] BL_UP[75] BL_UP[76] BL_UP[77] BL_UP[78] BL_UP[79]
+ BL_UP[80] BL_UP[81] BL_UP[82] BL_UP[83] BL_UP[84] BL_UP[85] BL_UP[86]
+ BL_UP[87] BL_UP[88] BL_UP[89] BL_UP[90] BL_UP[91] BL_UP[92] BL_UP[93]
+ BL_UP[94] BL_UP[95] BL_UP[96] BL_UP[97] BL_UP[98] BL_UP[99] BL_UP[100]
+ BL_UP[101] BL_UP[102] BL_UP[103] BL_UP[104] BL_UP[105] BL_UP[106] BL_UP[107]
+ BL_UP[108] BL_UP[109] BL_UP[110] BL_UP[111] BL_UP[112] BL_UP[113] BL_UP[114]
+ BL_UP[115] BL_UP[116] BL_UP[117] BL_UP[118] BL_UP[119] BL_UP[120] BL_UP[121]
+ BL_UP[122] BL_UP[123] BL_UP[124] BL_UP[125] BL_UP[126] BL_UP[127] BL_UP[128]
+ BL_UP[129] BL_UP[130] BL_UP[131] BL_UP[132] BL_UP[133] BL_UP[134] BL_UP[135]
+ BL_UP[136] BL_UP[137] BL_UP[138] BL_UP[139] BL_UP[140] BL_UP[141] BL_UP[142]
+ BL_UP[143] BL_UP[144] BL_UP[145] BL_UP[146] BL_UP[147] BL_UP[148] BL_UP[149]
+ BL_UP[150] BL_UP[151] BL_UP[152] BL_UP[153] BL_UP[154] BL_UP[155] BL_UP[156]
+ BL_UP[157] BL_UP[158] BL_UP[159] BL_UP[160] BL_UP[161] BL_UP[162] BL_UP[163]
+ BL_UP[164] BL_UP[165] BL_UP[166] BL_UP[167] BL_UP[168] BL_UP[169] BL_UP[170]
+ BL_UP[171] BL_UP[172] BL_UP[173] BL_UP[174] BL_UP[175] BL_UP[176] BL_UP[177]
+ BL_UP[178] BL_UP[179] BL_UP[180] BL_UP[181] BL_UP[182] BL_UP[183] BL_UP[184]
+ BL_UP[185] BL_UP[186] BL_UP[187] BL_UP[188] BL_UP[189] BL_UP[190] BL_UP[191]
+ BL_UP[192] BL_UP[193] BL_UP[194] BL_UP[195] BL_UP[196] BL_UP[197] BL_UP[198]
+ BL_UP[199] BL_UP[200] BL_UP[201] BL_UP[202] BL_UP[203] BL_UP[204] BL_UP[205]
+ BL_UP[206] BL_UP[207] BL_UP[208] BL_UP[209] BL_UP[210] BL_UP[211] BL_UP[212]
+ BL_UP[213] BL_UP[214] BL_UP[215] BL_UP[216] BL_UP[217] BL_UP[218] BL_UP[219]
+ BL_UP[220] BL_UP[221] BL_UP[222] BL_UP[223] BL_UP[224] BL_UP[225] BL_UP[226]
+ BL_UP[227] BL_UP[228] BL_UP[229] BL_UP[230] BL_UP[231] BL_UP[232] BL_UP[233]
+ BL_UP[234] BL_UP[235] BL_UP[236] BL_UP[237] BL_UP[238] BL_UP[239] BL_UP[240]
+ BL_UP[241] BL_UP[242] BL_UP[243] BL_UP[244] BL_UP[245] BL_UP[246] BL_UP[247]
+ BL_UP[248] BL_UP[249] BL_UP[250] BL_UP[251] BL_UP[252] BL_UP[253] BL_UP[254]
+ BL_UP[255] BL_UP[256] BL_UP[257] BL_UP[258] BL_UP[259] BL_UP[260] BL_UP[261]
+ BL_UP[262] BL_UP[263] BL_UP[264] BL_UP[265] BL_UP[266] BL_UP[267] BL_UP[268]
+ BL_UP[269] BL_UP[270] BL_UP[271] BL_UP[272] BL_UP[273] BL_UP[274] BL_UP[275]
+ BL_UP[276] BL_UP[277] BL_UP[278] BL_UP[279] BL_UP[280] BL_UP[281] BL_UP[282]
+ BL_UP[283] BL_UP[284] BL_UP[285] BL_UP[286] BL_UP[287] GBL[0] GBL[1] GBL[2]
+ GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12]
+ GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBLB[0] GBLB[1] GBLB[2] GBLB[3]
+ GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12]
+ GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9]
+ GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] LIOPD PDI PDOX
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
XLIO_M16_SD_0 BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5]
+ BLB_DN[6] BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12]
+ BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3]
+ BLB_UP[4] BLB_UP[5] BLB_UP[6] BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10]
+ BLB_UP[11] BLB_UP[12] BLB_UP[13] BLB_UP[14] BLB_UP[15] BLEQ_DN BLEQ_UP
+ BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7]
+ BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14] BL_DN[15]
+ BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] BL_UP[7]
+ BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14] BL_UP[15]
+ GBL[0] GBLB[0] GW[0] GWB[0] LIOPD LIOPD PDO0 PDO17 RE SAEB VXDDAI VDDI VSSI WE
+ YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6]
+ Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_1 BLB_DN[16] BLB_DN[17] BLB_DN[18] BLB_DN[19] BLB_DN[20] BLB_DN[21]
+ BLB_DN[22] BLB_DN[23] BLB_DN[24] BLB_DN[25] BLB_DN[26] BLB_DN[27] BLB_DN[28]
+ BLB_DN[29] BLB_DN[30] BLB_DN[31] BLB_UP[16] BLB_UP[17] BLB_UP[18] BLB_UP[19]
+ BLB_UP[20] BLB_UP[21] BLB_UP[22] BLB_UP[23] BLB_UP[24] BLB_UP[25] BLB_UP[26]
+ BLB_UP[27] BLB_UP[28] BLB_UP[29] BLB_UP[30] BLB_UP[31] BLEQ_DN BLEQ_UP
+ BL_DN[16] BL_DN[17] BL_DN[18] BL_DN[19] BL_DN[20] BL_DN[21] BL_DN[22]
+ BL_DN[23] BL_DN[24] BL_DN[25] BL_DN[26] BL_DN[27] BL_DN[28] BL_DN[29]
+ BL_DN[30] BL_DN[31] BL_UP[16] BL_UP[17] BL_UP[18] BL_UP[19] BL_UP[20]
+ BL_UP[21] BL_UP[22] BL_UP[23] BL_UP[24] BL_UP[25] BL_UP[26] BL_UP[27]
+ BL_UP[28] BL_UP[29] BL_UP[30] BL_UP[31] GBL[1] GBLB[1] GW[1] GWB[1] LIOPD PDO0
+ PDO1 PDO17 RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1]
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2]
+ Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_2 BLB_DN[32] BLB_DN[33] BLB_DN[34] BLB_DN[35] BLB_DN[36] BLB_DN[37]
+ BLB_DN[38] BLB_DN[39] BLB_DN[40] BLB_DN[41] BLB_DN[42] BLB_DN[43] BLB_DN[44]
+ BLB_DN[45] BLB_DN[46] BLB_DN[47] BLB_UP[32] BLB_UP[33] BLB_UP[34] BLB_UP[35]
+ BLB_UP[36] BLB_UP[37] BLB_UP[38] BLB_UP[39] BLB_UP[40] BLB_UP[41] BLB_UP[42]
+ BLB_UP[43] BLB_UP[44] BLB_UP[45] BLB_UP[46] BLB_UP[47] BLEQ_DN BLEQ_UP
+ BL_DN[32] BL_DN[33] BL_DN[34] BL_DN[35] BL_DN[36] BL_DN[37] BL_DN[38]
+ BL_DN[39] BL_DN[40] BL_DN[41] BL_DN[42] BL_DN[43] BL_DN[44] BL_DN[45]
+ BL_DN[46] BL_DN[47] BL_UP[32] BL_UP[33] BL_UP[34] BL_UP[35] BL_UP[36]
+ BL_UP[37] BL_UP[38] BL_UP[39] BL_UP[40] BL_UP[41] BL_UP[42] BL_UP[43]
+ BL_UP[44] BL_UP[45] BL_UP[46] BL_UP[47] GBL[2] GBLB[2] GW[2] GWB[2] LIOPD PDO1
+ PDO2 PDO17 RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1]
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2]
+ Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_3 BLB_DN[48] BLB_DN[49] BLB_DN[50] BLB_DN[51] BLB_DN[52] BLB_DN[53]
+ BLB_DN[54] BLB_DN[55] BLB_DN[56] BLB_DN[57] BLB_DN[58] BLB_DN[59] BLB_DN[60]
+ BLB_DN[61] BLB_DN[62] BLB_DN[63] BLB_UP[48] BLB_UP[49] BLB_UP[50] BLB_UP[51]
+ BLB_UP[52] BLB_UP[53] BLB_UP[54] BLB_UP[55] BLB_UP[56] BLB_UP[57] BLB_UP[58]
+ BLB_UP[59] BLB_UP[60] BLB_UP[61] BLB_UP[62] BLB_UP[63] BLEQ_DN BLEQ_UP
+ BL_DN[48] BL_DN[49] BL_DN[50] BL_DN[51] BL_DN[52] BL_DN[53] BL_DN[54]
+ BL_DN[55] BL_DN[56] BL_DN[57] BL_DN[58] BL_DN[59] BL_DN[60] BL_DN[61]
+ BL_DN[62] BL_DN[63] BL_UP[48] BL_UP[49] BL_UP[50] BL_UP[51] BL_UP[52]
+ BL_UP[53] BL_UP[54] BL_UP[55] BL_UP[56] BL_UP[57] BL_UP[58] BL_UP[59]
+ BL_UP[60] BL_UP[61] BL_UP[62] BL_UP[63] GBL[3] GBLB[3] GW[3] GWB[3] LIOPD PDO2
+ PDO3 PDO17 RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1]
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2]
+ Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_4 BLB_DN[64] BLB_DN[65] BLB_DN[66] BLB_DN[67] BLB_DN[68] BLB_DN[69]
+ BLB_DN[70] BLB_DN[71] BLB_DN[72] BLB_DN[73] BLB_DN[74] BLB_DN[75] BLB_DN[76]
+ BLB_DN[77] BLB_DN[78] BLB_DN[79] BLB_UP[64] BLB_UP[65] BLB_UP[66] BLB_UP[67]
+ BLB_UP[68] BLB_UP[69] BLB_UP[70] BLB_UP[71] BLB_UP[72] BLB_UP[73] BLB_UP[74]
+ BLB_UP[75] BLB_UP[76] BLB_UP[77] BLB_UP[78] BLB_UP[79] BLEQ_DN BLEQ_UP
+ BL_DN[64] BL_DN[65] BL_DN[66] BL_DN[67] BL_DN[68] BL_DN[69] BL_DN[70]
+ BL_DN[71] BL_DN[72] BL_DN[73] BL_DN[74] BL_DN[75] BL_DN[76] BL_DN[77]
+ BL_DN[78] BL_DN[79] BL_UP[64] BL_UP[65] BL_UP[66] BL_UP[67] BL_UP[68]
+ BL_UP[69] BL_UP[70] BL_UP[71] BL_UP[72] BL_UP[73] BL_UP[74] BL_UP[75]
+ BL_UP[76] BL_UP[77] BL_UP[78] BL_UP[79] GBL[4] GBLB[4] GW[4] GWB[4] LIOPD PDO3
+ PDO4 PDO17 RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1]
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2]
+ Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_5 BLB_DN[80] BLB_DN[81] BLB_DN[82] BLB_DN[83] BLB_DN[84] BLB_DN[85]
+ BLB_DN[86] BLB_DN[87] BLB_DN[88] BLB_DN[89] BLB_DN[90] BLB_DN[91] BLB_DN[92]
+ BLB_DN[93] BLB_DN[94] BLB_DN[95] BLB_UP[80] BLB_UP[81] BLB_UP[82] BLB_UP[83]
+ BLB_UP[84] BLB_UP[85] BLB_UP[86] BLB_UP[87] BLB_UP[88] BLB_UP[89] BLB_UP[90]
+ BLB_UP[91] BLB_UP[92] BLB_UP[93] BLB_UP[94] BLB_UP[95] BLEQ_DN BLEQ_UP
+ BL_DN[80] BL_DN[81] BL_DN[82] BL_DN[83] BL_DN[84] BL_DN[85] BL_DN[86]
+ BL_DN[87] BL_DN[88] BL_DN[89] BL_DN[90] BL_DN[91] BL_DN[92] BL_DN[93]
+ BL_DN[94] BL_DN[95] BL_UP[80] BL_UP[81] BL_UP[82] BL_UP[83] BL_UP[84]
+ BL_UP[85] BL_UP[86] BL_UP[87] BL_UP[88] BL_UP[89] BL_UP[90] BL_UP[91]
+ BL_UP[92] BL_UP[93] BL_UP[94] BL_UP[95] GBL[5] GBLB[5] GW[5] GWB[5] LIOPD PDO4
+ PDO5 PDO17 RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1]
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2]
+ Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_6 BLB_DN[96] BLB_DN[97] BLB_DN[98] BLB_DN[99] BLB_DN[100]
+ BLB_DN[101] BLB_DN[102] BLB_DN[103] BLB_DN[104] BLB_DN[105] BLB_DN[106]
+ BLB_DN[107] BLB_DN[108] BLB_DN[109] BLB_DN[110] BLB_DN[111] BLB_UP[96]
+ BLB_UP[97] BLB_UP[98] BLB_UP[99] BLB_UP[100] BLB_UP[101] BLB_UP[102]
+ BLB_UP[103] BLB_UP[104] BLB_UP[105] BLB_UP[106] BLB_UP[107] BLB_UP[108]
+ BLB_UP[109] BLB_UP[110] BLB_UP[111] BLEQ_DN BLEQ_UP BL_DN[96] BL_DN[97]
+ BL_DN[98] BL_DN[99] BL_DN[100] BL_DN[101] BL_DN[102] BL_DN[103] BL_DN[104]
+ BL_DN[105] BL_DN[106] BL_DN[107] BL_DN[108] BL_DN[109] BL_DN[110] BL_DN[111]
+ BL_UP[96] BL_UP[97] BL_UP[98] BL_UP[99] BL_UP[100] BL_UP[101] BL_UP[102]
+ BL_UP[103] BL_UP[104] BL_UP[105] BL_UP[106] BL_UP[107] BL_UP[108] BL_UP[109]
+ BL_UP[110] BL_UP[111] GBL[6] GBLB[6] GW[6] GWB[6] LIOPD PDO5 PDO6 PDO17 RE
+ SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_7 BLB_DN[112] BLB_DN[113] BLB_DN[114] BLB_DN[115] BLB_DN[116]
+ BLB_DN[117] BLB_DN[118] BLB_DN[119] BLB_DN[120] BLB_DN[121] BLB_DN[122]
+ BLB_DN[123] BLB_DN[124] BLB_DN[125] BLB_DN[126] BLB_DN[127] BLB_UP[112]
+ BLB_UP[113] BLB_UP[114] BLB_UP[115] BLB_UP[116] BLB_UP[117] BLB_UP[118]
+ BLB_UP[119] BLB_UP[120] BLB_UP[121] BLB_UP[122] BLB_UP[123] BLB_UP[124]
+ BLB_UP[125] BLB_UP[126] BLB_UP[127] BLEQ_DN BLEQ_UP BL_DN[112] BL_DN[113]
+ BL_DN[114] BL_DN[115] BL_DN[116] BL_DN[117] BL_DN[118] BL_DN[119] BL_DN[120]
+ BL_DN[121] BL_DN[122] BL_DN[123] BL_DN[124] BL_DN[125] BL_DN[126] BL_DN[127]
+ BL_UP[112] BL_UP[113] BL_UP[114] BL_UP[115] BL_UP[116] BL_UP[117] BL_UP[118]
+ BL_UP[119] BL_UP[120] BL_UP[121] BL_UP[122] BL_UP[123] BL_UP[124] BL_UP[125]
+ BL_UP[126] BL_UP[127] GBL[7] GBLB[7] GW[7] GWB[7] LIOPD PDO6 PDO7 PDO17 RE
+ SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_8 BLB_DN[128] BLB_DN[129] BLB_DN[130] BLB_DN[131] BLB_DN[132]
+ BLB_DN[133] BLB_DN[134] BLB_DN[135] BLB_DN[136] BLB_DN[137] BLB_DN[138]
+ BLB_DN[139] BLB_DN[140] BLB_DN[141] BLB_DN[142] BLB_DN[143] BLB_UP[128]
+ BLB_UP[129] BLB_UP[130] BLB_UP[131] BLB_UP[132] BLB_UP[133] BLB_UP[134]
+ BLB_UP[135] BLB_UP[136] BLB_UP[137] BLB_UP[138] BLB_UP[139] BLB_UP[140]
+ BLB_UP[141] BLB_UP[142] BLB_UP[143] BLEQ_DN BLEQ_UP BL_DN[128] BL_DN[129]
+ BL_DN[130] BL_DN[131] BL_DN[132] BL_DN[133] BL_DN[134] BL_DN[135] BL_DN[136]
+ BL_DN[137] BL_DN[138] BL_DN[139] BL_DN[140] BL_DN[141] BL_DN[142] BL_DN[143]
+ BL_UP[128] BL_UP[129] BL_UP[130] BL_UP[131] BL_UP[132] BL_UP[133] BL_UP[134]
+ BL_UP[135] BL_UP[136] BL_UP[137] BL_UP[138] BL_UP[139] BL_UP[140] BL_UP[141]
+ BL_UP[142] BL_UP[143] GBL[8] GBLB[8] GW[8] GWB[8] LIOPD PDO7 PDO8 PDO17 RE
+ SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_9 BLB_DN[144] BLB_DN[145] BLB_DN[146] BLB_DN[147] BLB_DN[148]
+ BLB_DN[149] BLB_DN[150] BLB_DN[151] BLB_DN[152] BLB_DN[153] BLB_DN[154]
+ BLB_DN[155] BLB_DN[156] BLB_DN[157] BLB_DN[158] BLB_DN[159] BLB_UP[144]
+ BLB_UP[145] BLB_UP[146] BLB_UP[147] BLB_UP[148] BLB_UP[149] BLB_UP[150]
+ BLB_UP[151] BLB_UP[152] BLB_UP[153] BLB_UP[154] BLB_UP[155] BLB_UP[156]
+ BLB_UP[157] BLB_UP[158] BLB_UP[159] BLEQ_DN BLEQ_UP BL_DN[144] BL_DN[145]
+ BL_DN[146] BL_DN[147] BL_DN[148] BL_DN[149] BL_DN[150] BL_DN[151] BL_DN[152]
+ BL_DN[153] BL_DN[154] BL_DN[155] BL_DN[156] BL_DN[157] BL_DN[158] BL_DN[159]
+ BL_UP[144] BL_UP[145] BL_UP[146] BL_UP[147] BL_UP[148] BL_UP[149] BL_UP[150]
+ BL_UP[151] BL_UP[152] BL_UP[153] BL_UP[154] BL_UP[155] BL_UP[156] BL_UP[157]
+ BL_UP[158] BL_UP[159] GBL[9] GBLB[9] GW[9] GWB[9] LIOPD PDO8 PDO9 PDO17 RE
+ SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_10 BLB_DN[160] BLB_DN[161] BLB_DN[162] BLB_DN[163] BLB_DN[164]
+ BLB_DN[165] BLB_DN[166] BLB_DN[167] BLB_DN[168] BLB_DN[169] BLB_DN[170]
+ BLB_DN[171] BLB_DN[172] BLB_DN[173] BLB_DN[174] BLB_DN[175] BLB_UP[160]
+ BLB_UP[161] BLB_UP[162] BLB_UP[163] BLB_UP[164] BLB_UP[165] BLB_UP[166]
+ BLB_UP[167] BLB_UP[168] BLB_UP[169] BLB_UP[170] BLB_UP[171] BLB_UP[172]
+ BLB_UP[173] BLB_UP[174] BLB_UP[175] BLEQ_DN BLEQ_UP BL_DN[160] BL_DN[161]
+ BL_DN[162] BL_DN[163] BL_DN[164] BL_DN[165] BL_DN[166] BL_DN[167] BL_DN[168]
+ BL_DN[169] BL_DN[170] BL_DN[171] BL_DN[172] BL_DN[173] BL_DN[174] BL_DN[175]
+ BL_UP[160] BL_UP[161] BL_UP[162] BL_UP[163] BL_UP[164] BL_UP[165] BL_UP[166]
+ BL_UP[167] BL_UP[168] BL_UP[169] BL_UP[170] BL_UP[171] BL_UP[172] BL_UP[173]
+ BL_UP[174] BL_UP[175] GBL[10] GBLB[10] GW[10] GWB[10] LIOPD PDO9 PDO10 PDO17
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_11 BLB_DN[176] BLB_DN[177] BLB_DN[178] BLB_DN[179] BLB_DN[180]
+ BLB_DN[181] BLB_DN[182] BLB_DN[183] BLB_DN[184] BLB_DN[185] BLB_DN[186]
+ BLB_DN[187] BLB_DN[188] BLB_DN[189] BLB_DN[190] BLB_DN[191] BLB_UP[176]
+ BLB_UP[177] BLB_UP[178] BLB_UP[179] BLB_UP[180] BLB_UP[181] BLB_UP[182]
+ BLB_UP[183] BLB_UP[184] BLB_UP[185] BLB_UP[186] BLB_UP[187] BLB_UP[188]
+ BLB_UP[189] BLB_UP[190] BLB_UP[191] BLEQ_DN BLEQ_UP BL_DN[176] BL_DN[177]
+ BL_DN[178] BL_DN[179] BL_DN[180] BL_DN[181] BL_DN[182] BL_DN[183] BL_DN[184]
+ BL_DN[185] BL_DN[186] BL_DN[187] BL_DN[188] BL_DN[189] BL_DN[190] BL_DN[191]
+ BL_UP[176] BL_UP[177] BL_UP[178] BL_UP[179] BL_UP[180] BL_UP[181] BL_UP[182]
+ BL_UP[183] BL_UP[184] BL_UP[185] BL_UP[186] BL_UP[187] BL_UP[188] BL_UP[189]
+ BL_UP[190] BL_UP[191] GBL[11] GBLB[11] GW[11] GWB[11] LIOPD PDO10 PDO11 PDO17
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_12 BLB_DN[192] BLB_DN[193] BLB_DN[194] BLB_DN[195] BLB_DN[196]
+ BLB_DN[197] BLB_DN[198] BLB_DN[199] BLB_DN[200] BLB_DN[201] BLB_DN[202]
+ BLB_DN[203] BLB_DN[204] BLB_DN[205] BLB_DN[206] BLB_DN[207] BLB_UP[192]
+ BLB_UP[193] BLB_UP[194] BLB_UP[195] BLB_UP[196] BLB_UP[197] BLB_UP[198]
+ BLB_UP[199] BLB_UP[200] BLB_UP[201] BLB_UP[202] BLB_UP[203] BLB_UP[204]
+ BLB_UP[205] BLB_UP[206] BLB_UP[207] BLEQ_DN BLEQ_UP BL_DN[192] BL_DN[193]
+ BL_DN[194] BL_DN[195] BL_DN[196] BL_DN[197] BL_DN[198] BL_DN[199] BL_DN[200]
+ BL_DN[201] BL_DN[202] BL_DN[203] BL_DN[204] BL_DN[205] BL_DN[206] BL_DN[207]
+ BL_UP[192] BL_UP[193] BL_UP[194] BL_UP[195] BL_UP[196] BL_UP[197] BL_UP[198]
+ BL_UP[199] BL_UP[200] BL_UP[201] BL_UP[202] BL_UP[203] BL_UP[204] BL_UP[205]
+ BL_UP[206] BL_UP[207] GBL[12] GBLB[12] GW[12] GWB[12] LIOPD PDO11 PDO12 PDO17
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_13 BLB_DN[208] BLB_DN[209] BLB_DN[210] BLB_DN[211] BLB_DN[212]
+ BLB_DN[213] BLB_DN[214] BLB_DN[215] BLB_DN[216] BLB_DN[217] BLB_DN[218]
+ BLB_DN[219] BLB_DN[220] BLB_DN[221] BLB_DN[222] BLB_DN[223] BLB_UP[208]
+ BLB_UP[209] BLB_UP[210] BLB_UP[211] BLB_UP[212] BLB_UP[213] BLB_UP[214]
+ BLB_UP[215] BLB_UP[216] BLB_UP[217] BLB_UP[218] BLB_UP[219] BLB_UP[220]
+ BLB_UP[221] BLB_UP[222] BLB_UP[223] BLEQ_DN BLEQ_UP BL_DN[208] BL_DN[209]
+ BL_DN[210] BL_DN[211] BL_DN[212] BL_DN[213] BL_DN[214] BL_DN[215] BL_DN[216]
+ BL_DN[217] BL_DN[218] BL_DN[219] BL_DN[220] BL_DN[221] BL_DN[222] BL_DN[223]
+ BL_UP[208] BL_UP[209] BL_UP[210] BL_UP[211] BL_UP[212] BL_UP[213] BL_UP[214]
+ BL_UP[215] BL_UP[216] BL_UP[217] BL_UP[218] BL_UP[219] BL_UP[220] BL_UP[221]
+ BL_UP[222] BL_UP[223] GBL[13] GBLB[13] GW[13] GWB[13] LIOPD PDO12 PDO13 PDO17
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_14 BLB_DN[224] BLB_DN[225] BLB_DN[226] BLB_DN[227] BLB_DN[228]
+ BLB_DN[229] BLB_DN[230] BLB_DN[231] BLB_DN[232] BLB_DN[233] BLB_DN[234]
+ BLB_DN[235] BLB_DN[236] BLB_DN[237] BLB_DN[238] BLB_DN[239] BLB_UP[224]
+ BLB_UP[225] BLB_UP[226] BLB_UP[227] BLB_UP[228] BLB_UP[229] BLB_UP[230]
+ BLB_UP[231] BLB_UP[232] BLB_UP[233] BLB_UP[234] BLB_UP[235] BLB_UP[236]
+ BLB_UP[237] BLB_UP[238] BLB_UP[239] BLEQ_DN BLEQ_UP BL_DN[224] BL_DN[225]
+ BL_DN[226] BL_DN[227] BL_DN[228] BL_DN[229] BL_DN[230] BL_DN[231] BL_DN[232]
+ BL_DN[233] BL_DN[234] BL_DN[235] BL_DN[236] BL_DN[237] BL_DN[238] BL_DN[239]
+ BL_UP[224] BL_UP[225] BL_UP[226] BL_UP[227] BL_UP[228] BL_UP[229] BL_UP[230]
+ BL_UP[231] BL_UP[232] BL_UP[233] BL_UP[234] BL_UP[235] BL_UP[236] BL_UP[237]
+ BL_UP[238] BL_UP[239] GBL[14] GBLB[14] GW[14] GWB[14] LIOPD PDO13 PDO14 PDO17
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_15 BLB_DN[240] BLB_DN[241] BLB_DN[242] BLB_DN[243] BLB_DN[244]
+ BLB_DN[245] BLB_DN[246] BLB_DN[247] BLB_DN[248] BLB_DN[249] BLB_DN[250]
+ BLB_DN[251] BLB_DN[252] BLB_DN[253] BLB_DN[254] BLB_DN[255] BLB_UP[240]
+ BLB_UP[241] BLB_UP[242] BLB_UP[243] BLB_UP[244] BLB_UP[245] BLB_UP[246]
+ BLB_UP[247] BLB_UP[248] BLB_UP[249] BLB_UP[250] BLB_UP[251] BLB_UP[252]
+ BLB_UP[253] BLB_UP[254] BLB_UP[255] BLEQ_DN BLEQ_UP BL_DN[240] BL_DN[241]
+ BL_DN[242] BL_DN[243] BL_DN[244] BL_DN[245] BL_DN[246] BL_DN[247] BL_DN[248]
+ BL_DN[249] BL_DN[250] BL_DN[251] BL_DN[252] BL_DN[253] BL_DN[254] BL_DN[255]
+ BL_UP[240] BL_UP[241] BL_UP[242] BL_UP[243] BL_UP[244] BL_UP[245] BL_UP[246]
+ BL_UP[247] BL_UP[248] BL_UP[249] BL_UP[250] BL_UP[251] BL_UP[252] BL_UP[253]
+ BL_UP[254] BL_UP[255] GBL[15] GBLB[15] GW[15] GWB[15] LIOPD PDO14 PDO15 PDO17
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_16 BLB_DN[256] BLB_DN[257] BLB_DN[258] BLB_DN[259] BLB_DN[260]
+ BLB_DN[261] BLB_DN[262] BLB_DN[263] BLB_DN[264] BLB_DN[265] BLB_DN[266]
+ BLB_DN[267] BLB_DN[268] BLB_DN[269] BLB_DN[270] BLB_DN[271] BLB_UP[256]
+ BLB_UP[257] BLB_UP[258] BLB_UP[259] BLB_UP[260] BLB_UP[261] BLB_UP[262]
+ BLB_UP[263] BLB_UP[264] BLB_UP[265] BLB_UP[266] BLB_UP[267] BLB_UP[268]
+ BLB_UP[269] BLB_UP[270] BLB_UP[271] BLEQ_DN BLEQ_UP BL_DN[256] BL_DN[257]
+ BL_DN[258] BL_DN[259] BL_DN[260] BL_DN[261] BL_DN[262] BL_DN[263] BL_DN[264]
+ BL_DN[265] BL_DN[266] BL_DN[267] BL_DN[268] BL_DN[269] BL_DN[270] BL_DN[271]
+ BL_UP[256] BL_UP[257] BL_UP[258] BL_UP[259] BL_UP[260] BL_UP[261] BL_UP[262]
+ BL_UP[263] BL_UP[264] BL_UP[265] BL_UP[266] BL_UP[267] BL_UP[268] BL_UP[269]
+ BL_UP[270] BL_UP[271] GBL[16] GBLB[16] GW[16] GWB[16] LIOPD PDO15 PDO16 PDO17
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
XLIO_M16_SD_17 BLB_DN[272] BLB_DN[273] BLB_DN[274] BLB_DN[275] BLB_DN[276]
+ BLB_DN[277] BLB_DN[278] BLB_DN[279] BLB_DN[280] BLB_DN[281] BLB_DN[282]
+ BLB_DN[283] BLB_DN[284] BLB_DN[285] BLB_DN[286] BLB_DN[287] BLB_UP[272]
+ BLB_UP[273] BLB_UP[274] BLB_UP[275] BLB_UP[276] BLB_UP[277] BLB_UP[278]
+ BLB_UP[279] BLB_UP[280] BLB_UP[281] BLB_UP[282] BLB_UP[283] BLB_UP[284]
+ BLB_UP[285] BLB_UP[286] BLB_UP[287] BLEQ_DN BLEQ_UP BL_DN[272] BL_DN[273]
+ BL_DN[274] BL_DN[275] BL_DN[276] BL_DN[277] BL_DN[278] BL_DN[279] BL_DN[280]
+ BL_DN[281] BL_DN[282] BL_DN[283] BL_DN[284] BL_DN[285] BL_DN[286] BL_DN[287]
+ BL_UP[272] BL_UP[273] BL_UP[274] BL_UP[275] BL_UP[276] BL_UP[277] BL_UP[278]
+ BL_UP[279] BL_UP[280] BL_UP[281] BL_UP[282] BL_UP[283] BL_UP[284] BL_UP[285]
+ BL_UP[286] BL_UP[287] GBL[17] GBLB[17] GW[17] GWB[17] LIOPD PDO16 PDO17 PDO17
+ RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1BSVTSWSO8000Y24_LIO_M16_SD
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_LIO_MCB_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6]
+ GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15]
+ GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23]
+ GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31]
+ GBLB[32] GBLB[33] GBLB[34] GBLB[35] VXDDAI LIOPD WL[0] WL[1] WL[2] WL[3] WL[4]
+ WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16]
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27]
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38]
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49]
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60]
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71]
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82]
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93]
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103]
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112]
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121]
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130]
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139]
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148]
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157]
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166]
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175]
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184]
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193]
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202]
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211]
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220]
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229]
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238]
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247]
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256]
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265]
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274]
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283]
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292]
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301]
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310]
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319]
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328]
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337]
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346]
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355]
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364]
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373]
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382]
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391]
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400]
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409]
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418]
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427]
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436]
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445]
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454]
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463]
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472]
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481]
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490]
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499]
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508]
+ WL[509] WL[510] WL[511] BLEQ_DN BLEQ_UP GW[0] GW[1] GW[2] GW[3] GW[4] GW[5]
+ GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2]
+ GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12]
+ GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21]
+ GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30]
+ GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] RE SAEB WE Y_DN[0] Y_DN[1] Y_DN[2]
+ Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3]
+ Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] YL_LIO[0] YL_LIO[1] VDDI VSSI
XCELL_ARR_DN_F BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6]
+ BL_DN[7] BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14]
+ BL_DN[15] BL_DN[16] BL_DN[17] BL_DN[18] BL_DN[19] BL_DN[20] BL_DN[21]
+ BL_DN[22] BL_DN[23] BL_DN[24] BL_DN[25] BL_DN[26] BL_DN[27] BL_DN[28]
+ BL_DN[29] BL_DN[30] BL_DN[31] BL_DN[32] BL_DN[33] BL_DN[34] BL_DN[35]
+ BL_DN[36] BL_DN[37] BL_DN[38] BL_DN[39] BL_DN[40] BL_DN[41] BL_DN[42]
+ BL_DN[43] BL_DN[44] BL_DN[45] BL_DN[46] BL_DN[47] BL_DN[48] BL_DN[49]
+ BL_DN[50] BL_DN[51] BL_DN[52] BL_DN[53] BL_DN[54] BL_DN[55] BL_DN[56]
+ BL_DN[57] BL_DN[58] BL_DN[59] BL_DN[60] BL_DN[61] BL_DN[62] BL_DN[63]
+ BL_DN[64] BL_DN[65] BL_DN[66] BL_DN[67] BL_DN[68] BL_DN[69] BL_DN[70]
+ BL_DN[71] BL_DN[72] BL_DN[73] BL_DN[74] BL_DN[75] BL_DN[76] BL_DN[77]
+ BL_DN[78] BL_DN[79] BL_DN[80] BL_DN[81] BL_DN[82] BL_DN[83] BL_DN[84]
+ BL_DN[85] BL_DN[86] BL_DN[87] BL_DN[88] BL_DN[89] BL_DN[90] BL_DN[91]
+ BL_DN[92] BL_DN[93] BL_DN[94] BL_DN[95] BL_DN[96] BL_DN[97] BL_DN[98]
+ BL_DN[99] BL_DN[100] BL_DN[101] BL_DN[102] BL_DN[103] BL_DN[104] BL_DN[105]
+ BL_DN[106] BL_DN[107] BL_DN[108] BL_DN[109] BL_DN[110] BL_DN[111] BL_DN[112]
+ BL_DN[113] BL_DN[114] BL_DN[115] BL_DN[116] BL_DN[117] BL_DN[118] BL_DN[119]
+ BL_DN[120] BL_DN[121] BL_DN[122] BL_DN[123] BL_DN[124] BL_DN[125] BL_DN[126]
+ BL_DN[127] BL_DN[128] BL_DN[129] BL_DN[130] BL_DN[131] BL_DN[132] BL_DN[133]
+ BL_DN[134] BL_DN[135] BL_DN[136] BL_DN[137] BL_DN[138] BL_DN[139] BL_DN[140]
+ BL_DN[141] BL_DN[142] BL_DN[143] BL_DN[144] BL_DN[145] BL_DN[146] BL_DN[147]
+ BL_DN[148] BL_DN[149] BL_DN[150] BL_DN[151] BL_DN[152] BL_DN[153] BL_DN[154]
+ BL_DN[155] BL_DN[156] BL_DN[157] BL_DN[158] BL_DN[159] BL_DN[160] BL_DN[161]
+ BL_DN[162] BL_DN[163] BL_DN[164] BL_DN[165] BL_DN[166] BL_DN[167] BL_DN[168]
+ BL_DN[169] BL_DN[170] BL_DN[171] BL_DN[172] BL_DN[173] BL_DN[174] BL_DN[175]
+ BL_DN[176] BL_DN[177] BL_DN[178] BL_DN[179] BL_DN[180] BL_DN[181] BL_DN[182]
+ BL_DN[183] BL_DN[184] BL_DN[185] BL_DN[186] BL_DN[187] BL_DN[188] BL_DN[189]
+ BL_DN[190] BL_DN[191] BL_DN[192] BL_DN[193] BL_DN[194] BL_DN[195] BL_DN[196]
+ BL_DN[197] BL_DN[198] BL_DN[199] BL_DN[200] BL_DN[201] BL_DN[202] BL_DN[203]
+ BL_DN[204] BL_DN[205] BL_DN[206] BL_DN[207] BL_DN[208] BL_DN[209] BL_DN[210]
+ BL_DN[211] BL_DN[212] BL_DN[213] BL_DN[214] BL_DN[215] BL_DN[216] BL_DN[217]
+ BL_DN[218] BL_DN[219] BL_DN[220] BL_DN[221] BL_DN[222] BL_DN[223] BL_DN[224]
+ BL_DN[225] BL_DN[226] BL_DN[227] BL_DN[228] BL_DN[229] BL_DN[230] BL_DN[231]
+ BL_DN[232] BL_DN[233] BL_DN[234] BL_DN[235] BL_DN[236] BL_DN[237] BL_DN[238]
+ BL_DN[239] BL_DN[240] BL_DN[241] BL_DN[242] BL_DN[243] BL_DN[244] BL_DN[245]
+ BL_DN[246] BL_DN[247] BL_DN[248] BL_DN[249] BL_DN[250] BL_DN[251] BL_DN[252]
+ BL_DN[253] BL_DN[254] BL_DN[255] BL_DN[256] BL_DN[257] BL_DN[258] BL_DN[259]
+ BL_DN[260] BL_DN[261] BL_DN[262] BL_DN[263] BL_DN[264] BL_DN[265] BL_DN[266]
+ BL_DN[267] BL_DN[268] BL_DN[269] BL_DN[270] BL_DN[271] BL_DN[272] BL_DN[273]
+ BL_DN[274] BL_DN[275] BL_DN[276] BL_DN[277] BL_DN[278] BL_DN[279] BL_DN[280]
+ BL_DN[281] BL_DN[282] BL_DN[283] BL_DN[284] BL_DN[285] BL_DN[286] BL_DN[287]
+ BL_DN[288] BL_DN[289] BL_DN[290] BL_DN[291] BL_DN[292] BL_DN[293] BL_DN[294]
+ BL_DN[295] BL_DN[296] BL_DN[297] BL_DN[298] BL_DN[299] BL_DN[300] BL_DN[301]
+ BL_DN[302] BL_DN[303] BL_DN[304] BL_DN[305] BL_DN[306] BL_DN[307] BL_DN[308]
+ BL_DN[309] BL_DN[310] BL_DN[311] BL_DN[312] BL_DN[313] BL_DN[314] BL_DN[315]
+ BL_DN[316] BL_DN[317] BL_DN[318] BL_DN[319] BL_DN[320] BL_DN[321] BL_DN[322]
+ BL_DN[323] BL_DN[324] BL_DN[325] BL_DN[326] BL_DN[327] BL_DN[328] BL_DN[329]
+ BL_DN[330] BL_DN[331] BL_DN[332] BL_DN[333] BL_DN[334] BL_DN[335] BL_DN[336]
+ BL_DN[337] BL_DN[338] BL_DN[339] BL_DN[340] BL_DN[341] BL_DN[342] BL_DN[343]
+ BL_DN[344] BL_DN[345] BL_DN[346] BL_DN[347] BL_DN[348] BL_DN[349] BL_DN[350]
+ BL_DN[351] BL_DN[352] BL_DN[353] BL_DN[354] BL_DN[355] BL_DN[356] BL_DN[357]
+ BL_DN[358] BL_DN[359] BL_DN[360] BL_DN[361] BL_DN[362] BL_DN[363] BL_DN[364]
+ BL_DN[365] BL_DN[366] BL_DN[367] BL_DN[368] BL_DN[369] BL_DN[370] BL_DN[371]
+ BL_DN[372] BL_DN[373] BL_DN[374] BL_DN[375] BL_DN[376] BL_DN[377] BL_DN[378]
+ BL_DN[379] BL_DN[380] BL_DN[381] BL_DN[382] BL_DN[383] BL_DN[384] BL_DN[385]
+ BL_DN[386] BL_DN[387] BL_DN[388] BL_DN[389] BL_DN[390] BL_DN[391] BL_DN[392]
+ BL_DN[393] BL_DN[394] BL_DN[395] BL_DN[396] BL_DN[397] BL_DN[398] BL_DN[399]
+ BL_DN[400] BL_DN[401] BL_DN[402] BL_DN[403] BL_DN[404] BL_DN[405] BL_DN[406]
+ BL_DN[407] BL_DN[408] BL_DN[409] BL_DN[410] BL_DN[411] BL_DN[412] BL_DN[413]
+ BL_DN[414] BL_DN[415] BL_DN[416] BL_DN[417] BL_DN[418] BL_DN[419] BL_DN[420]
+ BL_DN[421] BL_DN[422] BL_DN[423] BL_DN[424] BL_DN[425] BL_DN[426] BL_DN[427]
+ BL_DN[428] BL_DN[429] BL_DN[430] BL_DN[431] BL_DN[432] BL_DN[433] BL_DN[434]
+ BL_DN[435] BL_DN[436] BL_DN[437] BL_DN[438] BL_DN[439] BL_DN[440] BL_DN[441]
+ BL_DN[442] BL_DN[443] BL_DN[444] BL_DN[445] BL_DN[446] BL_DN[447] BL_DN[448]
+ BL_DN[449] BL_DN[450] BL_DN[451] BL_DN[452] BL_DN[453] BL_DN[454] BL_DN[455]
+ BL_DN[456] BL_DN[457] BL_DN[458] BL_DN[459] BL_DN[460] BL_DN[461] BL_DN[462]
+ BL_DN[463] BL_DN[464] BL_DN[465] BL_DN[466] BL_DN[467] BL_DN[468] BL_DN[469]
+ BL_DN[470] BL_DN[471] BL_DN[472] BL_DN[473] BL_DN[474] BL_DN[475] BL_DN[476]
+ BL_DN[477] BL_DN[478] BL_DN[479] BL_DN[480] BL_DN[481] BL_DN[482] BL_DN[483]
+ BL_DN[484] BL_DN[485] BL_DN[486] BL_DN[487] BL_DN[488] BL_DN[489] BL_DN[490]
+ BL_DN[491] BL_DN[492] BL_DN[493] BL_DN[494] BL_DN[495] BL_DN[496] BL_DN[497]
+ BL_DN[498] BL_DN[499] BL_DN[500] BL_DN[501] BL_DN[502] BL_DN[503] BL_DN[504]
+ BL_DN[505] BL_DN[506] BL_DN[507] BL_DN[508] BL_DN[509] BL_DN[510] BL_DN[511]
+ BL_DN[512] BL_DN[513] BL_DN[514] BL_DN[515] BL_DN[516] BL_DN[517] BL_DN[518]
+ BL_DN[519] BL_DN[520] BL_DN[521] BL_DN[522] BL_DN[523] BL_DN[524] BL_DN[525]
+ BL_DN[526] BL_DN[527] BL_DN[528] BL_DN[529] BL_DN[530] BL_DN[531] BL_DN[532]
+ BL_DN[533] BL_DN[534] BL_DN[535] BL_DN[536] BL_DN[537] BL_DN[538] BL_DN[539]
+ BL_DN[540] BL_DN[541] BL_DN[542] BL_DN[543] BL_DN[544] BL_DN[545] BL_DN[546]
+ BL_DN[547] BL_DN[548] BL_DN[549] BL_DN[550] BL_DN[551] BL_DN[552] BL_DN[553]
+ BL_DN[554] BL_DN[555] BL_DN[556] BL_DN[557] BL_DN[558] BL_DN[559] BL_DN[560]
+ BL_DN[561] BL_DN[562] BL_DN[563] BL_DN[564] BL_DN[565] BL_DN[566] BL_DN[567]
+ BL_DN[568] BL_DN[569] BL_DN[570] BL_DN[571] BL_DN[572] BL_DN[573] BL_DN[574]
+ BL_DN[575] BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5]
+ BLB_DN[6] BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12]
+ BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_DN[16] BLB_DN[17] BLB_DN[18] BLB_DN[19]
+ BLB_DN[20] BLB_DN[21] BLB_DN[22] BLB_DN[23] BLB_DN[24] BLB_DN[25] BLB_DN[26]
+ BLB_DN[27] BLB_DN[28] BLB_DN[29] BLB_DN[30] BLB_DN[31] BLB_DN[32] BLB_DN[33]
+ BLB_DN[34] BLB_DN[35] BLB_DN[36] BLB_DN[37] BLB_DN[38] BLB_DN[39] BLB_DN[40]
+ BLB_DN[41] BLB_DN[42] BLB_DN[43] BLB_DN[44] BLB_DN[45] BLB_DN[46] BLB_DN[47]
+ BLB_DN[48] BLB_DN[49] BLB_DN[50] BLB_DN[51] BLB_DN[52] BLB_DN[53] BLB_DN[54]
+ BLB_DN[55] BLB_DN[56] BLB_DN[57] BLB_DN[58] BLB_DN[59] BLB_DN[60] BLB_DN[61]
+ BLB_DN[62] BLB_DN[63] BLB_DN[64] BLB_DN[65] BLB_DN[66] BLB_DN[67] BLB_DN[68]
+ BLB_DN[69] BLB_DN[70] BLB_DN[71] BLB_DN[72] BLB_DN[73] BLB_DN[74] BLB_DN[75]
+ BLB_DN[76] BLB_DN[77] BLB_DN[78] BLB_DN[79] BLB_DN[80] BLB_DN[81] BLB_DN[82]
+ BLB_DN[83] BLB_DN[84] BLB_DN[85] BLB_DN[86] BLB_DN[87] BLB_DN[88] BLB_DN[89]
+ BLB_DN[90] BLB_DN[91] BLB_DN[92] BLB_DN[93] BLB_DN[94] BLB_DN[95] BLB_DN[96]
+ BLB_DN[97] BLB_DN[98] BLB_DN[99] BLB_DN[100] BLB_DN[101] BLB_DN[102]
+ BLB_DN[103] BLB_DN[104] BLB_DN[105] BLB_DN[106] BLB_DN[107] BLB_DN[108]
+ BLB_DN[109] BLB_DN[110] BLB_DN[111] BLB_DN[112] BLB_DN[113] BLB_DN[114]
+ BLB_DN[115] BLB_DN[116] BLB_DN[117] BLB_DN[118] BLB_DN[119] BLB_DN[120]
+ BLB_DN[121] BLB_DN[122] BLB_DN[123] BLB_DN[124] BLB_DN[125] BLB_DN[126]
+ BLB_DN[127] BLB_DN[128] BLB_DN[129] BLB_DN[130] BLB_DN[131] BLB_DN[132]
+ BLB_DN[133] BLB_DN[134] BLB_DN[135] BLB_DN[136] BLB_DN[137] BLB_DN[138]
+ BLB_DN[139] BLB_DN[140] BLB_DN[141] BLB_DN[142] BLB_DN[143] BLB_DN[144]
+ BLB_DN[145] BLB_DN[146] BLB_DN[147] BLB_DN[148] BLB_DN[149] BLB_DN[150]
+ BLB_DN[151] BLB_DN[152] BLB_DN[153] BLB_DN[154] BLB_DN[155] BLB_DN[156]
+ BLB_DN[157] BLB_DN[158] BLB_DN[159] BLB_DN[160] BLB_DN[161] BLB_DN[162]
+ BLB_DN[163] BLB_DN[164] BLB_DN[165] BLB_DN[166] BLB_DN[167] BLB_DN[168]
+ BLB_DN[169] BLB_DN[170] BLB_DN[171] BLB_DN[172] BLB_DN[173] BLB_DN[174]
+ BLB_DN[175] BLB_DN[176] BLB_DN[177] BLB_DN[178] BLB_DN[179] BLB_DN[180]
+ BLB_DN[181] BLB_DN[182] BLB_DN[183] BLB_DN[184] BLB_DN[185] BLB_DN[186]
+ BLB_DN[187] BLB_DN[188] BLB_DN[189] BLB_DN[190] BLB_DN[191] BLB_DN[192]
+ BLB_DN[193] BLB_DN[194] BLB_DN[195] BLB_DN[196] BLB_DN[197] BLB_DN[198]
+ BLB_DN[199] BLB_DN[200] BLB_DN[201] BLB_DN[202] BLB_DN[203] BLB_DN[204]
+ BLB_DN[205] BLB_DN[206] BLB_DN[207] BLB_DN[208] BLB_DN[209] BLB_DN[210]
+ BLB_DN[211] BLB_DN[212] BLB_DN[213] BLB_DN[214] BLB_DN[215] BLB_DN[216]
+ BLB_DN[217] BLB_DN[218] BLB_DN[219] BLB_DN[220] BLB_DN[221] BLB_DN[222]
+ BLB_DN[223] BLB_DN[224] BLB_DN[225] BLB_DN[226] BLB_DN[227] BLB_DN[228]
+ BLB_DN[229] BLB_DN[230] BLB_DN[231] BLB_DN[232] BLB_DN[233] BLB_DN[234]
+ BLB_DN[235] BLB_DN[236] BLB_DN[237] BLB_DN[238] BLB_DN[239] BLB_DN[240]
+ BLB_DN[241] BLB_DN[242] BLB_DN[243] BLB_DN[244] BLB_DN[245] BLB_DN[246]
+ BLB_DN[247] BLB_DN[248] BLB_DN[249] BLB_DN[250] BLB_DN[251] BLB_DN[252]
+ BLB_DN[253] BLB_DN[254] BLB_DN[255] BLB_DN[256] BLB_DN[257] BLB_DN[258]
+ BLB_DN[259] BLB_DN[260] BLB_DN[261] BLB_DN[262] BLB_DN[263] BLB_DN[264]
+ BLB_DN[265] BLB_DN[266] BLB_DN[267] BLB_DN[268] BLB_DN[269] BLB_DN[270]
+ BLB_DN[271] BLB_DN[272] BLB_DN[273] BLB_DN[274] BLB_DN[275] BLB_DN[276]
+ BLB_DN[277] BLB_DN[278] BLB_DN[279] BLB_DN[280] BLB_DN[281] BLB_DN[282]
+ BLB_DN[283] BLB_DN[284] BLB_DN[285] BLB_DN[286] BLB_DN[287] BLB_DN[288]
+ BLB_DN[289] BLB_DN[290] BLB_DN[291] BLB_DN[292] BLB_DN[293] BLB_DN[294]
+ BLB_DN[295] BLB_DN[296] BLB_DN[297] BLB_DN[298] BLB_DN[299] BLB_DN[300]
+ BLB_DN[301] BLB_DN[302] BLB_DN[303] BLB_DN[304] BLB_DN[305] BLB_DN[306]
+ BLB_DN[307] BLB_DN[308] BLB_DN[309] BLB_DN[310] BLB_DN[311] BLB_DN[312]
+ BLB_DN[313] BLB_DN[314] BLB_DN[315] BLB_DN[316] BLB_DN[317] BLB_DN[318]
+ BLB_DN[319] BLB_DN[320] BLB_DN[321] BLB_DN[322] BLB_DN[323] BLB_DN[324]
+ BLB_DN[325] BLB_DN[326] BLB_DN[327] BLB_DN[328] BLB_DN[329] BLB_DN[330]
+ BLB_DN[331] BLB_DN[332] BLB_DN[333] BLB_DN[334] BLB_DN[335] BLB_DN[336]
+ BLB_DN[337] BLB_DN[338] BLB_DN[339] BLB_DN[340] BLB_DN[341] BLB_DN[342]
+ BLB_DN[343] BLB_DN[344] BLB_DN[345] BLB_DN[346] BLB_DN[347] BLB_DN[348]
+ BLB_DN[349] BLB_DN[350] BLB_DN[351] BLB_DN[352] BLB_DN[353] BLB_DN[354]
+ BLB_DN[355] BLB_DN[356] BLB_DN[357] BLB_DN[358] BLB_DN[359] BLB_DN[360]
+ BLB_DN[361] BLB_DN[362] BLB_DN[363] BLB_DN[364] BLB_DN[365] BLB_DN[366]
+ BLB_DN[367] BLB_DN[368] BLB_DN[369] BLB_DN[370] BLB_DN[371] BLB_DN[372]
+ BLB_DN[373] BLB_DN[374] BLB_DN[375] BLB_DN[376] BLB_DN[377] BLB_DN[378]
+ BLB_DN[379] BLB_DN[380] BLB_DN[381] BLB_DN[382] BLB_DN[383] BLB_DN[384]
+ BLB_DN[385] BLB_DN[386] BLB_DN[387] BLB_DN[388] BLB_DN[389] BLB_DN[390]
+ BLB_DN[391] BLB_DN[392] BLB_DN[393] BLB_DN[394] BLB_DN[395] BLB_DN[396]
+ BLB_DN[397] BLB_DN[398] BLB_DN[399] BLB_DN[400] BLB_DN[401] BLB_DN[402]
+ BLB_DN[403] BLB_DN[404] BLB_DN[405] BLB_DN[406] BLB_DN[407] BLB_DN[408]
+ BLB_DN[409] BLB_DN[410] BLB_DN[411] BLB_DN[412] BLB_DN[413] BLB_DN[414]
+ BLB_DN[415] BLB_DN[416] BLB_DN[417] BLB_DN[418] BLB_DN[419] BLB_DN[420]
+ BLB_DN[421] BLB_DN[422] BLB_DN[423] BLB_DN[424] BLB_DN[425] BLB_DN[426]
+ BLB_DN[427] BLB_DN[428] BLB_DN[429] BLB_DN[430] BLB_DN[431] BLB_DN[432]
+ BLB_DN[433] BLB_DN[434] BLB_DN[435] BLB_DN[436] BLB_DN[437] BLB_DN[438]
+ BLB_DN[439] BLB_DN[440] BLB_DN[441] BLB_DN[442] BLB_DN[443] BLB_DN[444]
+ BLB_DN[445] BLB_DN[446] BLB_DN[447] BLB_DN[448] BLB_DN[449] BLB_DN[450]
+ BLB_DN[451] BLB_DN[452] BLB_DN[453] BLB_DN[454] BLB_DN[455] BLB_DN[456]
+ BLB_DN[457] BLB_DN[458] BLB_DN[459] BLB_DN[460] BLB_DN[461] BLB_DN[462]
+ BLB_DN[463] BLB_DN[464] BLB_DN[465] BLB_DN[466] BLB_DN[467] BLB_DN[468]
+ BLB_DN[469] BLB_DN[470] BLB_DN[471] BLB_DN[472] BLB_DN[473] BLB_DN[474]
+ BLB_DN[475] BLB_DN[476] BLB_DN[477] BLB_DN[478] BLB_DN[479] BLB_DN[480]
+ BLB_DN[481] BLB_DN[482] BLB_DN[483] BLB_DN[484] BLB_DN[485] BLB_DN[486]
+ BLB_DN[487] BLB_DN[488] BLB_DN[489] BLB_DN[490] BLB_DN[491] BLB_DN[492]
+ BLB_DN[493] BLB_DN[494] BLB_DN[495] BLB_DN[496] BLB_DN[497] BLB_DN[498]
+ BLB_DN[499] BLB_DN[500] BLB_DN[501] BLB_DN[502] BLB_DN[503] BLB_DN[504]
+ BLB_DN[505] BLB_DN[506] BLB_DN[507] BLB_DN[508] BLB_DN[509] BLB_DN[510]
+ BLB_DN[511] BLB_DN[512] BLB_DN[513] BLB_DN[514] BLB_DN[515] BLB_DN[516]
+ BLB_DN[517] BLB_DN[518] BLB_DN[519] BLB_DN[520] BLB_DN[521] BLB_DN[522]
+ BLB_DN[523] BLB_DN[524] BLB_DN[525] BLB_DN[526] BLB_DN[527] BLB_DN[528]
+ BLB_DN[529] BLB_DN[530] BLB_DN[531] BLB_DN[532] BLB_DN[533] BLB_DN[534]
+ BLB_DN[535] BLB_DN[536] BLB_DN[537] BLB_DN[538] BLB_DN[539] BLB_DN[540]
+ BLB_DN[541] BLB_DN[542] BLB_DN[543] BLB_DN[544] BLB_DN[545] BLB_DN[546]
+ BLB_DN[547] BLB_DN[548] BLB_DN[549] BLB_DN[550] BLB_DN[551] BLB_DN[552]
+ BLB_DN[553] BLB_DN[554] BLB_DN[555] BLB_DN[556] BLB_DN[557] BLB_DN[558]
+ BLB_DN[559] BLB_DN[560] BLB_DN[561] BLB_DN[562] BLB_DN[563] BLB_DN[564]
+ BLB_DN[565] BLB_DN[566] BLB_DN[567] BLB_DN[568] BLB_DN[569] BLB_DN[570]
+ BLB_DN[571] BLB_DN[572] BLB_DN[573] BLB_DN[574] BLB_DN[575] WL[0] WL[1] WL[2]
+ WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14]
+ WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25]
+ WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36]
+ WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47]
+ WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58]
+ WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69]
+ WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80]
+ WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91]
+ WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101]
+ WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110]
+ WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119]
+ WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128]
+ WL[129] WL[130] WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137]
+ WL[138] WL[139] WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146]
+ WL[147] WL[148] WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155]
+ WL[156] WL[157] WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164]
+ WL[165] WL[166] WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173]
+ WL[174] WL[175] WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182]
+ WL[183] WL[184] WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191]
+ WL[192] WL[193] WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200]
+ WL[201] WL[202] WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209]
+ WL[210] WL[211] WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218]
+ WL[219] WL[220] WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227]
+ WL[228] WL[229] WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236]
+ WL[237] WL[238] WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245]
+ WL[246] WL[247] WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254]
+ WL[255] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6]
+ GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16]
+ GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25]
+ GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34]
+ GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7]
+ GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16]
+ GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24]
+ GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32]
+ GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7]
+ GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18]
+ GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29]
+ GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4]
+ GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14]
+ GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23]
+ GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32]
+ GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_XY_F
XCELL_ARR_UP_F BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6]
+ BL_UP[7] BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14]
+ BL_UP[15] BL_UP[16] BL_UP[17] BL_UP[18] BL_UP[19] BL_UP[20] BL_UP[21]
+ BL_UP[22] BL_UP[23] BL_UP[24] BL_UP[25] BL_UP[26] BL_UP[27] BL_UP[28]
+ BL_UP[29] BL_UP[30] BL_UP[31] BL_UP[32] BL_UP[33] BL_UP[34] BL_UP[35]
+ BL_UP[36] BL_UP[37] BL_UP[38] BL_UP[39] BL_UP[40] BL_UP[41] BL_UP[42]
+ BL_UP[43] BL_UP[44] BL_UP[45] BL_UP[46] BL_UP[47] BL_UP[48] BL_UP[49]
+ BL_UP[50] BL_UP[51] BL_UP[52] BL_UP[53] BL_UP[54] BL_UP[55] BL_UP[56]
+ BL_UP[57] BL_UP[58] BL_UP[59] BL_UP[60] BL_UP[61] BL_UP[62] BL_UP[63]
+ BL_UP[64] BL_UP[65] BL_UP[66] BL_UP[67] BL_UP[68] BL_UP[69] BL_UP[70]
+ BL_UP[71] BL_UP[72] BL_UP[73] BL_UP[74] BL_UP[75] BL_UP[76] BL_UP[77]
+ BL_UP[78] BL_UP[79] BL_UP[80] BL_UP[81] BL_UP[82] BL_UP[83] BL_UP[84]
+ BL_UP[85] BL_UP[86] BL_UP[87] BL_UP[88] BL_UP[89] BL_UP[90] BL_UP[91]
+ BL_UP[92] BL_UP[93] BL_UP[94] BL_UP[95] BL_UP[96] BL_UP[97] BL_UP[98]
+ BL_UP[99] BL_UP[100] BL_UP[101] BL_UP[102] BL_UP[103] BL_UP[104] BL_UP[105]
+ BL_UP[106] BL_UP[107] BL_UP[108] BL_UP[109] BL_UP[110] BL_UP[111] BL_UP[112]
+ BL_UP[113] BL_UP[114] BL_UP[115] BL_UP[116] BL_UP[117] BL_UP[118] BL_UP[119]
+ BL_UP[120] BL_UP[121] BL_UP[122] BL_UP[123] BL_UP[124] BL_UP[125] BL_UP[126]
+ BL_UP[127] BL_UP[128] BL_UP[129] BL_UP[130] BL_UP[131] BL_UP[132] BL_UP[133]
+ BL_UP[134] BL_UP[135] BL_UP[136] BL_UP[137] BL_UP[138] BL_UP[139] BL_UP[140]
+ BL_UP[141] BL_UP[142] BL_UP[143] BL_UP[144] BL_UP[145] BL_UP[146] BL_UP[147]
+ BL_UP[148] BL_UP[149] BL_UP[150] BL_UP[151] BL_UP[152] BL_UP[153] BL_UP[154]
+ BL_UP[155] BL_UP[156] BL_UP[157] BL_UP[158] BL_UP[159] BL_UP[160] BL_UP[161]
+ BL_UP[162] BL_UP[163] BL_UP[164] BL_UP[165] BL_UP[166] BL_UP[167] BL_UP[168]
+ BL_UP[169] BL_UP[170] BL_UP[171] BL_UP[172] BL_UP[173] BL_UP[174] BL_UP[175]
+ BL_UP[176] BL_UP[177] BL_UP[178] BL_UP[179] BL_UP[180] BL_UP[181] BL_UP[182]
+ BL_UP[183] BL_UP[184] BL_UP[185] BL_UP[186] BL_UP[187] BL_UP[188] BL_UP[189]
+ BL_UP[190] BL_UP[191] BL_UP[192] BL_UP[193] BL_UP[194] BL_UP[195] BL_UP[196]
+ BL_UP[197] BL_UP[198] BL_UP[199] BL_UP[200] BL_UP[201] BL_UP[202] BL_UP[203]
+ BL_UP[204] BL_UP[205] BL_UP[206] BL_UP[207] BL_UP[208] BL_UP[209] BL_UP[210]
+ BL_UP[211] BL_UP[212] BL_UP[213] BL_UP[214] BL_UP[215] BL_UP[216] BL_UP[217]
+ BL_UP[218] BL_UP[219] BL_UP[220] BL_UP[221] BL_UP[222] BL_UP[223] BL_UP[224]
+ BL_UP[225] BL_UP[226] BL_UP[227] BL_UP[228] BL_UP[229] BL_UP[230] BL_UP[231]
+ BL_UP[232] BL_UP[233] BL_UP[234] BL_UP[235] BL_UP[236] BL_UP[237] BL_UP[238]
+ BL_UP[239] BL_UP[240] BL_UP[241] BL_UP[242] BL_UP[243] BL_UP[244] BL_UP[245]
+ BL_UP[246] BL_UP[247] BL_UP[248] BL_UP[249] BL_UP[250] BL_UP[251] BL_UP[252]
+ BL_UP[253] BL_UP[254] BL_UP[255] BL_UP[256] BL_UP[257] BL_UP[258] BL_UP[259]
+ BL_UP[260] BL_UP[261] BL_UP[262] BL_UP[263] BL_UP[264] BL_UP[265] BL_UP[266]
+ BL_UP[267] BL_UP[268] BL_UP[269] BL_UP[270] BL_UP[271] BL_UP[272] BL_UP[273]
+ BL_UP[274] BL_UP[275] BL_UP[276] BL_UP[277] BL_UP[278] BL_UP[279] BL_UP[280]
+ BL_UP[281] BL_UP[282] BL_UP[283] BL_UP[284] BL_UP[285] BL_UP[286] BL_UP[287]
+ BL_UP[288] BL_UP[289] BL_UP[290] BL_UP[291] BL_UP[292] BL_UP[293] BL_UP[294]
+ BL_UP[295] BL_UP[296] BL_UP[297] BL_UP[298] BL_UP[299] BL_UP[300] BL_UP[301]
+ BL_UP[302] BL_UP[303] BL_UP[304] BL_UP[305] BL_UP[306] BL_UP[307] BL_UP[308]
+ BL_UP[309] BL_UP[310] BL_UP[311] BL_UP[312] BL_UP[313] BL_UP[314] BL_UP[315]
+ BL_UP[316] BL_UP[317] BL_UP[318] BL_UP[319] BL_UP[320] BL_UP[321] BL_UP[322]
+ BL_UP[323] BL_UP[324] BL_UP[325] BL_UP[326] BL_UP[327] BL_UP[328] BL_UP[329]
+ BL_UP[330] BL_UP[331] BL_UP[332] BL_UP[333] BL_UP[334] BL_UP[335] BL_UP[336]
+ BL_UP[337] BL_UP[338] BL_UP[339] BL_UP[340] BL_UP[341] BL_UP[342] BL_UP[343]
+ BL_UP[344] BL_UP[345] BL_UP[346] BL_UP[347] BL_UP[348] BL_UP[349] BL_UP[350]
+ BL_UP[351] BL_UP[352] BL_UP[353] BL_UP[354] BL_UP[355] BL_UP[356] BL_UP[357]
+ BL_UP[358] BL_UP[359] BL_UP[360] BL_UP[361] BL_UP[362] BL_UP[363] BL_UP[364]
+ BL_UP[365] BL_UP[366] BL_UP[367] BL_UP[368] BL_UP[369] BL_UP[370] BL_UP[371]
+ BL_UP[372] BL_UP[373] BL_UP[374] BL_UP[375] BL_UP[376] BL_UP[377] BL_UP[378]
+ BL_UP[379] BL_UP[380] BL_UP[381] BL_UP[382] BL_UP[383] BL_UP[384] BL_UP[385]
+ BL_UP[386] BL_UP[387] BL_UP[388] BL_UP[389] BL_UP[390] BL_UP[391] BL_UP[392]
+ BL_UP[393] BL_UP[394] BL_UP[395] BL_UP[396] BL_UP[397] BL_UP[398] BL_UP[399]
+ BL_UP[400] BL_UP[401] BL_UP[402] BL_UP[403] BL_UP[404] BL_UP[405] BL_UP[406]
+ BL_UP[407] BL_UP[408] BL_UP[409] BL_UP[410] BL_UP[411] BL_UP[412] BL_UP[413]
+ BL_UP[414] BL_UP[415] BL_UP[416] BL_UP[417] BL_UP[418] BL_UP[419] BL_UP[420]
+ BL_UP[421] BL_UP[422] BL_UP[423] BL_UP[424] BL_UP[425] BL_UP[426] BL_UP[427]
+ BL_UP[428] BL_UP[429] BL_UP[430] BL_UP[431] BL_UP[432] BL_UP[433] BL_UP[434]
+ BL_UP[435] BL_UP[436] BL_UP[437] BL_UP[438] BL_UP[439] BL_UP[440] BL_UP[441]
+ BL_UP[442] BL_UP[443] BL_UP[444] BL_UP[445] BL_UP[446] BL_UP[447] BL_UP[448]
+ BL_UP[449] BL_UP[450] BL_UP[451] BL_UP[452] BL_UP[453] BL_UP[454] BL_UP[455]
+ BL_UP[456] BL_UP[457] BL_UP[458] BL_UP[459] BL_UP[460] BL_UP[461] BL_UP[462]
+ BL_UP[463] BL_UP[464] BL_UP[465] BL_UP[466] BL_UP[467] BL_UP[468] BL_UP[469]
+ BL_UP[470] BL_UP[471] BL_UP[472] BL_UP[473] BL_UP[474] BL_UP[475] BL_UP[476]
+ BL_UP[477] BL_UP[478] BL_UP[479] BL_UP[480] BL_UP[481] BL_UP[482] BL_UP[483]
+ BL_UP[484] BL_UP[485] BL_UP[486] BL_UP[487] BL_UP[488] BL_UP[489] BL_UP[490]
+ BL_UP[491] BL_UP[492] BL_UP[493] BL_UP[494] BL_UP[495] BL_UP[496] BL_UP[497]
+ BL_UP[498] BL_UP[499] BL_UP[500] BL_UP[501] BL_UP[502] BL_UP[503] BL_UP[504]
+ BL_UP[505] BL_UP[506] BL_UP[507] BL_UP[508] BL_UP[509] BL_UP[510] BL_UP[511]
+ BL_UP[512] BL_UP[513] BL_UP[514] BL_UP[515] BL_UP[516] BL_UP[517] BL_UP[518]
+ BL_UP[519] BL_UP[520] BL_UP[521] BL_UP[522] BL_UP[523] BL_UP[524] BL_UP[525]
+ BL_UP[526] BL_UP[527] BL_UP[528] BL_UP[529] BL_UP[530] BL_UP[531] BL_UP[532]
+ BL_UP[533] BL_UP[534] BL_UP[535] BL_UP[536] BL_UP[537] BL_UP[538] BL_UP[539]
+ BL_UP[540] BL_UP[541] BL_UP[542] BL_UP[543] BL_UP[544] BL_UP[545] BL_UP[546]
+ BL_UP[547] BL_UP[548] BL_UP[549] BL_UP[550] BL_UP[551] BL_UP[552] BL_UP[553]
+ BL_UP[554] BL_UP[555] BL_UP[556] BL_UP[557] BL_UP[558] BL_UP[559] BL_UP[560]
+ BL_UP[561] BL_UP[562] BL_UP[563] BL_UP[564] BL_UP[565] BL_UP[566] BL_UP[567]
+ BL_UP[568] BL_UP[569] BL_UP[570] BL_UP[571] BL_UP[572] BL_UP[573] BL_UP[574]
+ BL_UP[575] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] BLB_UP[4] BLB_UP[5]
+ BLB_UP[6] BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10] BLB_UP[11] BLB_UP[12]
+ BLB_UP[13] BLB_UP[14] BLB_UP[15] BLB_UP[16] BLB_UP[17] BLB_UP[18] BLB_UP[19]
+ BLB_UP[20] BLB_UP[21] BLB_UP[22] BLB_UP[23] BLB_UP[24] BLB_UP[25] BLB_UP[26]
+ BLB_UP[27] BLB_UP[28] BLB_UP[29] BLB_UP[30] BLB_UP[31] BLB_UP[32] BLB_UP[33]
+ BLB_UP[34] BLB_UP[35] BLB_UP[36] BLB_UP[37] BLB_UP[38] BLB_UP[39] BLB_UP[40]
+ BLB_UP[41] BLB_UP[42] BLB_UP[43] BLB_UP[44] BLB_UP[45] BLB_UP[46] BLB_UP[47]
+ BLB_UP[48] BLB_UP[49] BLB_UP[50] BLB_UP[51] BLB_UP[52] BLB_UP[53] BLB_UP[54]
+ BLB_UP[55] BLB_UP[56] BLB_UP[57] BLB_UP[58] BLB_UP[59] BLB_UP[60] BLB_UP[61]
+ BLB_UP[62] BLB_UP[63] BLB_UP[64] BLB_UP[65] BLB_UP[66] BLB_UP[67] BLB_UP[68]
+ BLB_UP[69] BLB_UP[70] BLB_UP[71] BLB_UP[72] BLB_UP[73] BLB_UP[74] BLB_UP[75]
+ BLB_UP[76] BLB_UP[77] BLB_UP[78] BLB_UP[79] BLB_UP[80] BLB_UP[81] BLB_UP[82]
+ BLB_UP[83] BLB_UP[84] BLB_UP[85] BLB_UP[86] BLB_UP[87] BLB_UP[88] BLB_UP[89]
+ BLB_UP[90] BLB_UP[91] BLB_UP[92] BLB_UP[93] BLB_UP[94] BLB_UP[95] BLB_UP[96]
+ BLB_UP[97] BLB_UP[98] BLB_UP[99] BLB_UP[100] BLB_UP[101] BLB_UP[102]
+ BLB_UP[103] BLB_UP[104] BLB_UP[105] BLB_UP[106] BLB_UP[107] BLB_UP[108]
+ BLB_UP[109] BLB_UP[110] BLB_UP[111] BLB_UP[112] BLB_UP[113] BLB_UP[114]
+ BLB_UP[115] BLB_UP[116] BLB_UP[117] BLB_UP[118] BLB_UP[119] BLB_UP[120]
+ BLB_UP[121] BLB_UP[122] BLB_UP[123] BLB_UP[124] BLB_UP[125] BLB_UP[126]
+ BLB_UP[127] BLB_UP[128] BLB_UP[129] BLB_UP[130] BLB_UP[131] BLB_UP[132]
+ BLB_UP[133] BLB_UP[134] BLB_UP[135] BLB_UP[136] BLB_UP[137] BLB_UP[138]
+ BLB_UP[139] BLB_UP[140] BLB_UP[141] BLB_UP[142] BLB_UP[143] BLB_UP[144]
+ BLB_UP[145] BLB_UP[146] BLB_UP[147] BLB_UP[148] BLB_UP[149] BLB_UP[150]
+ BLB_UP[151] BLB_UP[152] BLB_UP[153] BLB_UP[154] BLB_UP[155] BLB_UP[156]
+ BLB_UP[157] BLB_UP[158] BLB_UP[159] BLB_UP[160] BLB_UP[161] BLB_UP[162]
+ BLB_UP[163] BLB_UP[164] BLB_UP[165] BLB_UP[166] BLB_UP[167] BLB_UP[168]
+ BLB_UP[169] BLB_UP[170] BLB_UP[171] BLB_UP[172] BLB_UP[173] BLB_UP[174]
+ BLB_UP[175] BLB_UP[176] BLB_UP[177] BLB_UP[178] BLB_UP[179] BLB_UP[180]
+ BLB_UP[181] BLB_UP[182] BLB_UP[183] BLB_UP[184] BLB_UP[185] BLB_UP[186]
+ BLB_UP[187] BLB_UP[188] BLB_UP[189] BLB_UP[190] BLB_UP[191] BLB_UP[192]
+ BLB_UP[193] BLB_UP[194] BLB_UP[195] BLB_UP[196] BLB_UP[197] BLB_UP[198]
+ BLB_UP[199] BLB_UP[200] BLB_UP[201] BLB_UP[202] BLB_UP[203] BLB_UP[204]
+ BLB_UP[205] BLB_UP[206] BLB_UP[207] BLB_UP[208] BLB_UP[209] BLB_UP[210]
+ BLB_UP[211] BLB_UP[212] BLB_UP[213] BLB_UP[214] BLB_UP[215] BLB_UP[216]
+ BLB_UP[217] BLB_UP[218] BLB_UP[219] BLB_UP[220] BLB_UP[221] BLB_UP[222]
+ BLB_UP[223] BLB_UP[224] BLB_UP[225] BLB_UP[226] BLB_UP[227] BLB_UP[228]
+ BLB_UP[229] BLB_UP[230] BLB_UP[231] BLB_UP[232] BLB_UP[233] BLB_UP[234]
+ BLB_UP[235] BLB_UP[236] BLB_UP[237] BLB_UP[238] BLB_UP[239] BLB_UP[240]
+ BLB_UP[241] BLB_UP[242] BLB_UP[243] BLB_UP[244] BLB_UP[245] BLB_UP[246]
+ BLB_UP[247] BLB_UP[248] BLB_UP[249] BLB_UP[250] BLB_UP[251] BLB_UP[252]
+ BLB_UP[253] BLB_UP[254] BLB_UP[255] BLB_UP[256] BLB_UP[257] BLB_UP[258]
+ BLB_UP[259] BLB_UP[260] BLB_UP[261] BLB_UP[262] BLB_UP[263] BLB_UP[264]
+ BLB_UP[265] BLB_UP[266] BLB_UP[267] BLB_UP[268] BLB_UP[269] BLB_UP[270]
+ BLB_UP[271] BLB_UP[272] BLB_UP[273] BLB_UP[274] BLB_UP[275] BLB_UP[276]
+ BLB_UP[277] BLB_UP[278] BLB_UP[279] BLB_UP[280] BLB_UP[281] BLB_UP[282]
+ BLB_UP[283] BLB_UP[284] BLB_UP[285] BLB_UP[286] BLB_UP[287] BLB_UP[288]
+ BLB_UP[289] BLB_UP[290] BLB_UP[291] BLB_UP[292] BLB_UP[293] BLB_UP[294]
+ BLB_UP[295] BLB_UP[296] BLB_UP[297] BLB_UP[298] BLB_UP[299] BLB_UP[300]
+ BLB_UP[301] BLB_UP[302] BLB_UP[303] BLB_UP[304] BLB_UP[305] BLB_UP[306]
+ BLB_UP[307] BLB_UP[308] BLB_UP[309] BLB_UP[310] BLB_UP[311] BLB_UP[312]
+ BLB_UP[313] BLB_UP[314] BLB_UP[315] BLB_UP[316] BLB_UP[317] BLB_UP[318]
+ BLB_UP[319] BLB_UP[320] BLB_UP[321] BLB_UP[322] BLB_UP[323] BLB_UP[324]
+ BLB_UP[325] BLB_UP[326] BLB_UP[327] BLB_UP[328] BLB_UP[329] BLB_UP[330]
+ BLB_UP[331] BLB_UP[332] BLB_UP[333] BLB_UP[334] BLB_UP[335] BLB_UP[336]
+ BLB_UP[337] BLB_UP[338] BLB_UP[339] BLB_UP[340] BLB_UP[341] BLB_UP[342]
+ BLB_UP[343] BLB_UP[344] BLB_UP[345] BLB_UP[346] BLB_UP[347] BLB_UP[348]
+ BLB_UP[349] BLB_UP[350] BLB_UP[351] BLB_UP[352] BLB_UP[353] BLB_UP[354]
+ BLB_UP[355] BLB_UP[356] BLB_UP[357] BLB_UP[358] BLB_UP[359] BLB_UP[360]
+ BLB_UP[361] BLB_UP[362] BLB_UP[363] BLB_UP[364] BLB_UP[365] BLB_UP[366]
+ BLB_UP[367] BLB_UP[368] BLB_UP[369] BLB_UP[370] BLB_UP[371] BLB_UP[372]
+ BLB_UP[373] BLB_UP[374] BLB_UP[375] BLB_UP[376] BLB_UP[377] BLB_UP[378]
+ BLB_UP[379] BLB_UP[380] BLB_UP[381] BLB_UP[382] BLB_UP[383] BLB_UP[384]
+ BLB_UP[385] BLB_UP[386] BLB_UP[387] BLB_UP[388] BLB_UP[389] BLB_UP[390]
+ BLB_UP[391] BLB_UP[392] BLB_UP[393] BLB_UP[394] BLB_UP[395] BLB_UP[396]
+ BLB_UP[397] BLB_UP[398] BLB_UP[399] BLB_UP[400] BLB_UP[401] BLB_UP[402]
+ BLB_UP[403] BLB_UP[404] BLB_UP[405] BLB_UP[406] BLB_UP[407] BLB_UP[408]
+ BLB_UP[409] BLB_UP[410] BLB_UP[411] BLB_UP[412] BLB_UP[413] BLB_UP[414]
+ BLB_UP[415] BLB_UP[416] BLB_UP[417] BLB_UP[418] BLB_UP[419] BLB_UP[420]
+ BLB_UP[421] BLB_UP[422] BLB_UP[423] BLB_UP[424] BLB_UP[425] BLB_UP[426]
+ BLB_UP[427] BLB_UP[428] BLB_UP[429] BLB_UP[430] BLB_UP[431] BLB_UP[432]
+ BLB_UP[433] BLB_UP[434] BLB_UP[435] BLB_UP[436] BLB_UP[437] BLB_UP[438]
+ BLB_UP[439] BLB_UP[440] BLB_UP[441] BLB_UP[442] BLB_UP[443] BLB_UP[444]
+ BLB_UP[445] BLB_UP[446] BLB_UP[447] BLB_UP[448] BLB_UP[449] BLB_UP[450]
+ BLB_UP[451] BLB_UP[452] BLB_UP[453] BLB_UP[454] BLB_UP[455] BLB_UP[456]
+ BLB_UP[457] BLB_UP[458] BLB_UP[459] BLB_UP[460] BLB_UP[461] BLB_UP[462]
+ BLB_UP[463] BLB_UP[464] BLB_UP[465] BLB_UP[466] BLB_UP[467] BLB_UP[468]
+ BLB_UP[469] BLB_UP[470] BLB_UP[471] BLB_UP[472] BLB_UP[473] BLB_UP[474]
+ BLB_UP[475] BLB_UP[476] BLB_UP[477] BLB_UP[478] BLB_UP[479] BLB_UP[480]
+ BLB_UP[481] BLB_UP[482] BLB_UP[483] BLB_UP[484] BLB_UP[485] BLB_UP[486]
+ BLB_UP[487] BLB_UP[488] BLB_UP[489] BLB_UP[490] BLB_UP[491] BLB_UP[492]
+ BLB_UP[493] BLB_UP[494] BLB_UP[495] BLB_UP[496] BLB_UP[497] BLB_UP[498]
+ BLB_UP[499] BLB_UP[500] BLB_UP[501] BLB_UP[502] BLB_UP[503] BLB_UP[504]
+ BLB_UP[505] BLB_UP[506] BLB_UP[507] BLB_UP[508] BLB_UP[509] BLB_UP[510]
+ BLB_UP[511] BLB_UP[512] BLB_UP[513] BLB_UP[514] BLB_UP[515] BLB_UP[516]
+ BLB_UP[517] BLB_UP[518] BLB_UP[519] BLB_UP[520] BLB_UP[521] BLB_UP[522]
+ BLB_UP[523] BLB_UP[524] BLB_UP[525] BLB_UP[526] BLB_UP[527] BLB_UP[528]
+ BLB_UP[529] BLB_UP[530] BLB_UP[531] BLB_UP[532] BLB_UP[533] BLB_UP[534]
+ BLB_UP[535] BLB_UP[536] BLB_UP[537] BLB_UP[538] BLB_UP[539] BLB_UP[540]
+ BLB_UP[541] BLB_UP[542] BLB_UP[543] BLB_UP[544] BLB_UP[545] BLB_UP[546]
+ BLB_UP[547] BLB_UP[548] BLB_UP[549] BLB_UP[550] BLB_UP[551] BLB_UP[552]
+ BLB_UP[553] BLB_UP[554] BLB_UP[555] BLB_UP[556] BLB_UP[557] BLB_UP[558]
+ BLB_UP[559] BLB_UP[560] BLB_UP[561] BLB_UP[562] BLB_UP[563] BLB_UP[564]
+ BLB_UP[565] BLB_UP[566] BLB_UP[567] BLB_UP[568] BLB_UP[569] BLB_UP[570]
+ BLB_UP[571] BLB_UP[572] BLB_UP[573] BLB_UP[574] BLB_UP[575] WL[256] WL[257]
+ WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] WL[266]
+ WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] WL[275]
+ WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] WL[284]
+ WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] WL[293]
+ WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] WL[302]
+ WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] WL[311]
+ WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] WL[320]
+ WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] WL[329]
+ WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] WL[338]
+ WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] WL[347]
+ WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] WL[356]
+ WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] WL[365]
+ WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] WL[374]
+ WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] WL[383]
+ WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] WL[392]
+ WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] WL[401]
+ WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] WL[410]
+ WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] WL[419]
+ WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] WL[428]
+ WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] WL[437]
+ WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] WL[446]
+ WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] WL[455]
+ WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] WL[464]
+ WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] WL[473]
+ WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] WL[482]
+ WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] WL[491]
+ WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] WL[500]
+ WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] WL[509]
+ WL[510] WL[511] VXDDAI VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6]
+ GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15]
+ GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23]
+ GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31]
+ GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6]
+ GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17]
+ GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28]
+ GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3]
+ GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13]
+ GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22]
+ GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31]
+ GWB[32] GWB[33] GWB[34] GWB[35] S1BSVTSWSO8000Y24_CELL_ARR_XY_F
XLIO_L_SD BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] BLB_DN[6]
+ BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12] BLB_DN[13]
+ BLB_DN[14] BLB_DN[15] BLB_DN[16] BLB_DN[17] BLB_DN[18] BLB_DN[19] BLB_DN[20]
+ BLB_DN[21] BLB_DN[22] BLB_DN[23] BLB_DN[24] BLB_DN[25] BLB_DN[26] BLB_DN[27]
+ BLB_DN[28] BLB_DN[29] BLB_DN[30] BLB_DN[31] BLB_DN[32] BLB_DN[33] BLB_DN[34]
+ BLB_DN[35] BLB_DN[36] BLB_DN[37] BLB_DN[38] BLB_DN[39] BLB_DN[40] BLB_DN[41]
+ BLB_DN[42] BLB_DN[43] BLB_DN[44] BLB_DN[45] BLB_DN[46] BLB_DN[47] BLB_DN[48]
+ BLB_DN[49] BLB_DN[50] BLB_DN[51] BLB_DN[52] BLB_DN[53] BLB_DN[54] BLB_DN[55]
+ BLB_DN[56] BLB_DN[57] BLB_DN[58] BLB_DN[59] BLB_DN[60] BLB_DN[61] BLB_DN[62]
+ BLB_DN[63] BLB_DN[64] BLB_DN[65] BLB_DN[66] BLB_DN[67] BLB_DN[68] BLB_DN[69]
+ BLB_DN[70] BLB_DN[71] BLB_DN[72] BLB_DN[73] BLB_DN[74] BLB_DN[75] BLB_DN[76]
+ BLB_DN[77] BLB_DN[78] BLB_DN[79] BLB_DN[80] BLB_DN[81] BLB_DN[82] BLB_DN[83]
+ BLB_DN[84] BLB_DN[85] BLB_DN[86] BLB_DN[87] BLB_DN[88] BLB_DN[89] BLB_DN[90]
+ BLB_DN[91] BLB_DN[92] BLB_DN[93] BLB_DN[94] BLB_DN[95] BLB_DN[96] BLB_DN[97]
+ BLB_DN[98] BLB_DN[99] BLB_DN[100] BLB_DN[101] BLB_DN[102] BLB_DN[103]
+ BLB_DN[104] BLB_DN[105] BLB_DN[106] BLB_DN[107] BLB_DN[108] BLB_DN[109]
+ BLB_DN[110] BLB_DN[111] BLB_DN[112] BLB_DN[113] BLB_DN[114] BLB_DN[115]
+ BLB_DN[116] BLB_DN[117] BLB_DN[118] BLB_DN[119] BLB_DN[120] BLB_DN[121]
+ BLB_DN[122] BLB_DN[123] BLB_DN[124] BLB_DN[125] BLB_DN[126] BLB_DN[127]
+ BLB_DN[128] BLB_DN[129] BLB_DN[130] BLB_DN[131] BLB_DN[132] BLB_DN[133]
+ BLB_DN[134] BLB_DN[135] BLB_DN[136] BLB_DN[137] BLB_DN[138] BLB_DN[139]
+ BLB_DN[140] BLB_DN[141] BLB_DN[142] BLB_DN[143] BLB_DN[144] BLB_DN[145]
+ BLB_DN[146] BLB_DN[147] BLB_DN[148] BLB_DN[149] BLB_DN[150] BLB_DN[151]
+ BLB_DN[152] BLB_DN[153] BLB_DN[154] BLB_DN[155] BLB_DN[156] BLB_DN[157]
+ BLB_DN[158] BLB_DN[159] BLB_DN[160] BLB_DN[161] BLB_DN[162] BLB_DN[163]
+ BLB_DN[164] BLB_DN[165] BLB_DN[166] BLB_DN[167] BLB_DN[168] BLB_DN[169]
+ BLB_DN[170] BLB_DN[171] BLB_DN[172] BLB_DN[173] BLB_DN[174] BLB_DN[175]
+ BLB_DN[176] BLB_DN[177] BLB_DN[178] BLB_DN[179] BLB_DN[180] BLB_DN[181]
+ BLB_DN[182] BLB_DN[183] BLB_DN[184] BLB_DN[185] BLB_DN[186] BLB_DN[187]
+ BLB_DN[188] BLB_DN[189] BLB_DN[190] BLB_DN[191] BLB_DN[192] BLB_DN[193]
+ BLB_DN[194] BLB_DN[195] BLB_DN[196] BLB_DN[197] BLB_DN[198] BLB_DN[199]
+ BLB_DN[200] BLB_DN[201] BLB_DN[202] BLB_DN[203] BLB_DN[204] BLB_DN[205]
+ BLB_DN[206] BLB_DN[207] BLB_DN[208] BLB_DN[209] BLB_DN[210] BLB_DN[211]
+ BLB_DN[212] BLB_DN[213] BLB_DN[214] BLB_DN[215] BLB_DN[216] BLB_DN[217]
+ BLB_DN[218] BLB_DN[219] BLB_DN[220] BLB_DN[221] BLB_DN[222] BLB_DN[223]
+ BLB_DN[224] BLB_DN[225] BLB_DN[226] BLB_DN[227] BLB_DN[228] BLB_DN[229]
+ BLB_DN[230] BLB_DN[231] BLB_DN[232] BLB_DN[233] BLB_DN[234] BLB_DN[235]
+ BLB_DN[236] BLB_DN[237] BLB_DN[238] BLB_DN[239] BLB_DN[240] BLB_DN[241]
+ BLB_DN[242] BLB_DN[243] BLB_DN[244] BLB_DN[245] BLB_DN[246] BLB_DN[247]
+ BLB_DN[248] BLB_DN[249] BLB_DN[250] BLB_DN[251] BLB_DN[252] BLB_DN[253]
+ BLB_DN[254] BLB_DN[255] BLB_DN[256] BLB_DN[257] BLB_DN[258] BLB_DN[259]
+ BLB_DN[260] BLB_DN[261] BLB_DN[262] BLB_DN[263] BLB_DN[264] BLB_DN[265]
+ BLB_DN[266] BLB_DN[267] BLB_DN[268] BLB_DN[269] BLB_DN[270] BLB_DN[271]
+ BLB_DN[272] BLB_DN[273] BLB_DN[274] BLB_DN[275] BLB_DN[276] BLB_DN[277]
+ BLB_DN[278] BLB_DN[279] BLB_DN[280] BLB_DN[281] BLB_DN[282] BLB_DN[283]
+ BLB_DN[284] BLB_DN[285] BLB_DN[286] BLB_DN[287] BLB_UP[0] BLB_UP[1] BLB_UP[2]
+ BLB_UP[3] BLB_UP[4] BLB_UP[5] BLB_UP[6] BLB_UP[7] BLB_UP[8] BLB_UP[9]
+ BLB_UP[10] BLB_UP[11] BLB_UP[12] BLB_UP[13] BLB_UP[14] BLB_UP[15] BLB_UP[16]
+ BLB_UP[17] BLB_UP[18] BLB_UP[19] BLB_UP[20] BLB_UP[21] BLB_UP[22] BLB_UP[23]
+ BLB_UP[24] BLB_UP[25] BLB_UP[26] BLB_UP[27] BLB_UP[28] BLB_UP[29] BLB_UP[30]
+ BLB_UP[31] BLB_UP[32] BLB_UP[33] BLB_UP[34] BLB_UP[35] BLB_UP[36] BLB_UP[37]
+ BLB_UP[38] BLB_UP[39] BLB_UP[40] BLB_UP[41] BLB_UP[42] BLB_UP[43] BLB_UP[44]
+ BLB_UP[45] BLB_UP[46] BLB_UP[47] BLB_UP[48] BLB_UP[49] BLB_UP[50] BLB_UP[51]
+ BLB_UP[52] BLB_UP[53] BLB_UP[54] BLB_UP[55] BLB_UP[56] BLB_UP[57] BLB_UP[58]
+ BLB_UP[59] BLB_UP[60] BLB_UP[61] BLB_UP[62] BLB_UP[63] BLB_UP[64] BLB_UP[65]
+ BLB_UP[66] BLB_UP[67] BLB_UP[68] BLB_UP[69] BLB_UP[70] BLB_UP[71] BLB_UP[72]
+ BLB_UP[73] BLB_UP[74] BLB_UP[75] BLB_UP[76] BLB_UP[77] BLB_UP[78] BLB_UP[79]
+ BLB_UP[80] BLB_UP[81] BLB_UP[82] BLB_UP[83] BLB_UP[84] BLB_UP[85] BLB_UP[86]
+ BLB_UP[87] BLB_UP[88] BLB_UP[89] BLB_UP[90] BLB_UP[91] BLB_UP[92] BLB_UP[93]
+ BLB_UP[94] BLB_UP[95] BLB_UP[96] BLB_UP[97] BLB_UP[98] BLB_UP[99] BLB_UP[100]
+ BLB_UP[101] BLB_UP[102] BLB_UP[103] BLB_UP[104] BLB_UP[105] BLB_UP[106]
+ BLB_UP[107] BLB_UP[108] BLB_UP[109] BLB_UP[110] BLB_UP[111] BLB_UP[112]
+ BLB_UP[113] BLB_UP[114] BLB_UP[115] BLB_UP[116] BLB_UP[117] BLB_UP[118]
+ BLB_UP[119] BLB_UP[120] BLB_UP[121] BLB_UP[122] BLB_UP[123] BLB_UP[124]
+ BLB_UP[125] BLB_UP[126] BLB_UP[127] BLB_UP[128] BLB_UP[129] BLB_UP[130]
+ BLB_UP[131] BLB_UP[132] BLB_UP[133] BLB_UP[134] BLB_UP[135] BLB_UP[136]
+ BLB_UP[137] BLB_UP[138] BLB_UP[139] BLB_UP[140] BLB_UP[141] BLB_UP[142]
+ BLB_UP[143] BLB_UP[144] BLB_UP[145] BLB_UP[146] BLB_UP[147] BLB_UP[148]
+ BLB_UP[149] BLB_UP[150] BLB_UP[151] BLB_UP[152] BLB_UP[153] BLB_UP[154]
+ BLB_UP[155] BLB_UP[156] BLB_UP[157] BLB_UP[158] BLB_UP[159] BLB_UP[160]
+ BLB_UP[161] BLB_UP[162] BLB_UP[163] BLB_UP[164] BLB_UP[165] BLB_UP[166]
+ BLB_UP[167] BLB_UP[168] BLB_UP[169] BLB_UP[170] BLB_UP[171] BLB_UP[172]
+ BLB_UP[173] BLB_UP[174] BLB_UP[175] BLB_UP[176] BLB_UP[177] BLB_UP[178]
+ BLB_UP[179] BLB_UP[180] BLB_UP[181] BLB_UP[182] BLB_UP[183] BLB_UP[184]
+ BLB_UP[185] BLB_UP[186] BLB_UP[187] BLB_UP[188] BLB_UP[189] BLB_UP[190]
+ BLB_UP[191] BLB_UP[192] BLB_UP[193] BLB_UP[194] BLB_UP[195] BLB_UP[196]
+ BLB_UP[197] BLB_UP[198] BLB_UP[199] BLB_UP[200] BLB_UP[201] BLB_UP[202]
+ BLB_UP[203] BLB_UP[204] BLB_UP[205] BLB_UP[206] BLB_UP[207] BLB_UP[208]
+ BLB_UP[209] BLB_UP[210] BLB_UP[211] BLB_UP[212] BLB_UP[213] BLB_UP[214]
+ BLB_UP[215] BLB_UP[216] BLB_UP[217] BLB_UP[218] BLB_UP[219] BLB_UP[220]
+ BLB_UP[221] BLB_UP[222] BLB_UP[223] BLB_UP[224] BLB_UP[225] BLB_UP[226]
+ BLB_UP[227] BLB_UP[228] BLB_UP[229] BLB_UP[230] BLB_UP[231] BLB_UP[232]
+ BLB_UP[233] BLB_UP[234] BLB_UP[235] BLB_UP[236] BLB_UP[237] BLB_UP[238]
+ BLB_UP[239] BLB_UP[240] BLB_UP[241] BLB_UP[242] BLB_UP[243] BLB_UP[244]
+ BLB_UP[245] BLB_UP[246] BLB_UP[247] BLB_UP[248] BLB_UP[249] BLB_UP[250]
+ BLB_UP[251] BLB_UP[252] BLB_UP[253] BLB_UP[254] BLB_UP[255] BLB_UP[256]
+ BLB_UP[257] BLB_UP[258] BLB_UP[259] BLB_UP[260] BLB_UP[261] BLB_UP[262]
+ BLB_UP[263] BLB_UP[264] BLB_UP[265] BLB_UP[266] BLB_UP[267] BLB_UP[268]
+ BLB_UP[269] BLB_UP[270] BLB_UP[271] BLB_UP[272] BLB_UP[273] BLB_UP[274]
+ BLB_UP[275] BLB_UP[276] BLB_UP[277] BLB_UP[278] BLB_UP[279] BLB_UP[280]
+ BLB_UP[281] BLB_UP[282] BLB_UP[283] BLB_UP[284] BLB_UP[285] BLB_UP[286]
+ BLB_UP[287] BLEQ_DN BLEQ_UP BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4]
+ BL_DN[5] BL_DN[6] BL_DN[7] BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12]
+ BL_DN[13] BL_DN[14] BL_DN[15] BL_DN[16] BL_DN[17] BL_DN[18] BL_DN[19]
+ BL_DN[20] BL_DN[21] BL_DN[22] BL_DN[23] BL_DN[24] BL_DN[25] BL_DN[26]
+ BL_DN[27] BL_DN[28] BL_DN[29] BL_DN[30] BL_DN[31] BL_DN[32] BL_DN[33]
+ BL_DN[34] BL_DN[35] BL_DN[36] BL_DN[37] BL_DN[38] BL_DN[39] BL_DN[40]
+ BL_DN[41] BL_DN[42] BL_DN[43] BL_DN[44] BL_DN[45] BL_DN[46] BL_DN[47]
+ BL_DN[48] BL_DN[49] BL_DN[50] BL_DN[51] BL_DN[52] BL_DN[53] BL_DN[54]
+ BL_DN[55] BL_DN[56] BL_DN[57] BL_DN[58] BL_DN[59] BL_DN[60] BL_DN[61]
+ BL_DN[62] BL_DN[63] BL_DN[64] BL_DN[65] BL_DN[66] BL_DN[67] BL_DN[68]
+ BL_DN[69] BL_DN[70] BL_DN[71] BL_DN[72] BL_DN[73] BL_DN[74] BL_DN[75]
+ BL_DN[76] BL_DN[77] BL_DN[78] BL_DN[79] BL_DN[80] BL_DN[81] BL_DN[82]
+ BL_DN[83] BL_DN[84] BL_DN[85] BL_DN[86] BL_DN[87] BL_DN[88] BL_DN[89]
+ BL_DN[90] BL_DN[91] BL_DN[92] BL_DN[93] BL_DN[94] BL_DN[95] BL_DN[96]
+ BL_DN[97] BL_DN[98] BL_DN[99] BL_DN[100] BL_DN[101] BL_DN[102] BL_DN[103]
+ BL_DN[104] BL_DN[105] BL_DN[106] BL_DN[107] BL_DN[108] BL_DN[109] BL_DN[110]
+ BL_DN[111] BL_DN[112] BL_DN[113] BL_DN[114] BL_DN[115] BL_DN[116] BL_DN[117]
+ BL_DN[118] BL_DN[119] BL_DN[120] BL_DN[121] BL_DN[122] BL_DN[123] BL_DN[124]
+ BL_DN[125] BL_DN[126] BL_DN[127] BL_DN[128] BL_DN[129] BL_DN[130] BL_DN[131]
+ BL_DN[132] BL_DN[133] BL_DN[134] BL_DN[135] BL_DN[136] BL_DN[137] BL_DN[138]
+ BL_DN[139] BL_DN[140] BL_DN[141] BL_DN[142] BL_DN[143] BL_DN[144] BL_DN[145]
+ BL_DN[146] BL_DN[147] BL_DN[148] BL_DN[149] BL_DN[150] BL_DN[151] BL_DN[152]
+ BL_DN[153] BL_DN[154] BL_DN[155] BL_DN[156] BL_DN[157] BL_DN[158] BL_DN[159]
+ BL_DN[160] BL_DN[161] BL_DN[162] BL_DN[163] BL_DN[164] BL_DN[165] BL_DN[166]
+ BL_DN[167] BL_DN[168] BL_DN[169] BL_DN[170] BL_DN[171] BL_DN[172] BL_DN[173]
+ BL_DN[174] BL_DN[175] BL_DN[176] BL_DN[177] BL_DN[178] BL_DN[179] BL_DN[180]
+ BL_DN[181] BL_DN[182] BL_DN[183] BL_DN[184] BL_DN[185] BL_DN[186] BL_DN[187]
+ BL_DN[188] BL_DN[189] BL_DN[190] BL_DN[191] BL_DN[192] BL_DN[193] BL_DN[194]
+ BL_DN[195] BL_DN[196] BL_DN[197] BL_DN[198] BL_DN[199] BL_DN[200] BL_DN[201]
+ BL_DN[202] BL_DN[203] BL_DN[204] BL_DN[205] BL_DN[206] BL_DN[207] BL_DN[208]
+ BL_DN[209] BL_DN[210] BL_DN[211] BL_DN[212] BL_DN[213] BL_DN[214] BL_DN[215]
+ BL_DN[216] BL_DN[217] BL_DN[218] BL_DN[219] BL_DN[220] BL_DN[221] BL_DN[222]
+ BL_DN[223] BL_DN[224] BL_DN[225] BL_DN[226] BL_DN[227] BL_DN[228] BL_DN[229]
+ BL_DN[230] BL_DN[231] BL_DN[232] BL_DN[233] BL_DN[234] BL_DN[235] BL_DN[236]
+ BL_DN[237] BL_DN[238] BL_DN[239] BL_DN[240] BL_DN[241] BL_DN[242] BL_DN[243]
+ BL_DN[244] BL_DN[245] BL_DN[246] BL_DN[247] BL_DN[248] BL_DN[249] BL_DN[250]
+ BL_DN[251] BL_DN[252] BL_DN[253] BL_DN[254] BL_DN[255] BL_DN[256] BL_DN[257]
+ BL_DN[258] BL_DN[259] BL_DN[260] BL_DN[261] BL_DN[262] BL_DN[263] BL_DN[264]
+ BL_DN[265] BL_DN[266] BL_DN[267] BL_DN[268] BL_DN[269] BL_DN[270] BL_DN[271]
+ BL_DN[272] BL_DN[273] BL_DN[274] BL_DN[275] BL_DN[276] BL_DN[277] BL_DN[278]
+ BL_DN[279] BL_DN[280] BL_DN[281] BL_DN[282] BL_DN[283] BL_DN[284] BL_DN[285]
+ BL_DN[286] BL_DN[287] BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5]
+ BL_UP[6] BL_UP[7] BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13]
+ BL_UP[14] BL_UP[15] BL_UP[16] BL_UP[17] BL_UP[18] BL_UP[19] BL_UP[20]
+ BL_UP[21] BL_UP[22] BL_UP[23] BL_UP[24] BL_UP[25] BL_UP[26] BL_UP[27]
+ BL_UP[28] BL_UP[29] BL_UP[30] BL_UP[31] BL_UP[32] BL_UP[33] BL_UP[34]
+ BL_UP[35] BL_UP[36] BL_UP[37] BL_UP[38] BL_UP[39] BL_UP[40] BL_UP[41]
+ BL_UP[42] BL_UP[43] BL_UP[44] BL_UP[45] BL_UP[46] BL_UP[47] BL_UP[48]
+ BL_UP[49] BL_UP[50] BL_UP[51] BL_UP[52] BL_UP[53] BL_UP[54] BL_UP[55]
+ BL_UP[56] BL_UP[57] BL_UP[58] BL_UP[59] BL_UP[60] BL_UP[61] BL_UP[62]
+ BL_UP[63] BL_UP[64] BL_UP[65] BL_UP[66] BL_UP[67] BL_UP[68] BL_UP[69]
+ BL_UP[70] BL_UP[71] BL_UP[72] BL_UP[73] BL_UP[74] BL_UP[75] BL_UP[76]
+ BL_UP[77] BL_UP[78] BL_UP[79] BL_UP[80] BL_UP[81] BL_UP[82] BL_UP[83]
+ BL_UP[84] BL_UP[85] BL_UP[86] BL_UP[87] BL_UP[88] BL_UP[89] BL_UP[90]
+ BL_UP[91] BL_UP[92] BL_UP[93] BL_UP[94] BL_UP[95] BL_UP[96] BL_UP[97]
+ BL_UP[98] BL_UP[99] BL_UP[100] BL_UP[101] BL_UP[102] BL_UP[103] BL_UP[104]
+ BL_UP[105] BL_UP[106] BL_UP[107] BL_UP[108] BL_UP[109] BL_UP[110] BL_UP[111]
+ BL_UP[112] BL_UP[113] BL_UP[114] BL_UP[115] BL_UP[116] BL_UP[117] BL_UP[118]
+ BL_UP[119] BL_UP[120] BL_UP[121] BL_UP[122] BL_UP[123] BL_UP[124] BL_UP[125]
+ BL_UP[126] BL_UP[127] BL_UP[128] BL_UP[129] BL_UP[130] BL_UP[131] BL_UP[132]
+ BL_UP[133] BL_UP[134] BL_UP[135] BL_UP[136] BL_UP[137] BL_UP[138] BL_UP[139]
+ BL_UP[140] BL_UP[141] BL_UP[142] BL_UP[143] BL_UP[144] BL_UP[145] BL_UP[146]
+ BL_UP[147] BL_UP[148] BL_UP[149] BL_UP[150] BL_UP[151] BL_UP[152] BL_UP[153]
+ BL_UP[154] BL_UP[155] BL_UP[156] BL_UP[157] BL_UP[158] BL_UP[159] BL_UP[160]
+ BL_UP[161] BL_UP[162] BL_UP[163] BL_UP[164] BL_UP[165] BL_UP[166] BL_UP[167]
+ BL_UP[168] BL_UP[169] BL_UP[170] BL_UP[171] BL_UP[172] BL_UP[173] BL_UP[174]
+ BL_UP[175] BL_UP[176] BL_UP[177] BL_UP[178] BL_UP[179] BL_UP[180] BL_UP[181]
+ BL_UP[182] BL_UP[183] BL_UP[184] BL_UP[185] BL_UP[186] BL_UP[187] BL_UP[188]
+ BL_UP[189] BL_UP[190] BL_UP[191] BL_UP[192] BL_UP[193] BL_UP[194] BL_UP[195]
+ BL_UP[196] BL_UP[197] BL_UP[198] BL_UP[199] BL_UP[200] BL_UP[201] BL_UP[202]
+ BL_UP[203] BL_UP[204] BL_UP[205] BL_UP[206] BL_UP[207] BL_UP[208] BL_UP[209]
+ BL_UP[210] BL_UP[211] BL_UP[212] BL_UP[213] BL_UP[214] BL_UP[215] BL_UP[216]
+ BL_UP[217] BL_UP[218] BL_UP[219] BL_UP[220] BL_UP[221] BL_UP[222] BL_UP[223]
+ BL_UP[224] BL_UP[225] BL_UP[226] BL_UP[227] BL_UP[228] BL_UP[229] BL_UP[230]
+ BL_UP[231] BL_UP[232] BL_UP[233] BL_UP[234] BL_UP[235] BL_UP[236] BL_UP[237]
+ BL_UP[238] BL_UP[239] BL_UP[240] BL_UP[241] BL_UP[242] BL_UP[243] BL_UP[244]
+ BL_UP[245] BL_UP[246] BL_UP[247] BL_UP[248] BL_UP[249] BL_UP[250] BL_UP[251]
+ BL_UP[252] BL_UP[253] BL_UP[254] BL_UP[255] BL_UP[256] BL_UP[257] BL_UP[258]
+ BL_UP[259] BL_UP[260] BL_UP[261] BL_UP[262] BL_UP[263] BL_UP[264] BL_UP[265]
+ BL_UP[266] BL_UP[267] BL_UP[268] BL_UP[269] BL_UP[270] BL_UP[271] BL_UP[272]
+ BL_UP[273] BL_UP[274] BL_UP[275] BL_UP[276] BL_UP[277] BL_UP[278] BL_UP[279]
+ BL_UP[280] BL_UP[281] BL_UP[282] BL_UP[283] BL_UP[284] BL_UP[285] BL_UP[286]
+ BL_UP[287] GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8]
+ GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5]
+ GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15]
+ GWB[16] GWB[17] LIOPD LIOPD PDOXL RE SAEB VXDDAI VDDI VSSI WE YL_LIO[0]
+ YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7]
+ Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ S1BSVTSWSO8000Y24_LIO_L_SD
XLIO_R_SD BLB_DN[288] BLB_DN[289] BLB_DN[290] BLB_DN[291] BLB_DN[292]
+ BLB_DN[293] BLB_DN[294] BLB_DN[295] BLB_DN[296] BLB_DN[297] BLB_DN[298]
+ BLB_DN[299] BLB_DN[300] BLB_DN[301] BLB_DN[302] BLB_DN[303] BLB_DN[304]
+ BLB_DN[305] BLB_DN[306] BLB_DN[307] BLB_DN[308] BLB_DN[309] BLB_DN[310]
+ BLB_DN[311] BLB_DN[312] BLB_DN[313] BLB_DN[314] BLB_DN[315] BLB_DN[316]
+ BLB_DN[317] BLB_DN[318] BLB_DN[319] BLB_DN[320] BLB_DN[321] BLB_DN[322]
+ BLB_DN[323] BLB_DN[324] BLB_DN[325] BLB_DN[326] BLB_DN[327] BLB_DN[328]
+ BLB_DN[329] BLB_DN[330] BLB_DN[331] BLB_DN[332] BLB_DN[333] BLB_DN[334]
+ BLB_DN[335] BLB_DN[336] BLB_DN[337] BLB_DN[338] BLB_DN[339] BLB_DN[340]
+ BLB_DN[341] BLB_DN[342] BLB_DN[343] BLB_DN[344] BLB_DN[345] BLB_DN[346]
+ BLB_DN[347] BLB_DN[348] BLB_DN[349] BLB_DN[350] BLB_DN[351] BLB_DN[352]
+ BLB_DN[353] BLB_DN[354] BLB_DN[355] BLB_DN[356] BLB_DN[357] BLB_DN[358]
+ BLB_DN[359] BLB_DN[360] BLB_DN[361] BLB_DN[362] BLB_DN[363] BLB_DN[364]
+ BLB_DN[365] BLB_DN[366] BLB_DN[367] BLB_DN[368] BLB_DN[369] BLB_DN[370]
+ BLB_DN[371] BLB_DN[372] BLB_DN[373] BLB_DN[374] BLB_DN[375] BLB_DN[376]
+ BLB_DN[377] BLB_DN[378] BLB_DN[379] BLB_DN[380] BLB_DN[381] BLB_DN[382]
+ BLB_DN[383] BLB_DN[384] BLB_DN[385] BLB_DN[386] BLB_DN[387] BLB_DN[388]
+ BLB_DN[389] BLB_DN[390] BLB_DN[391] BLB_DN[392] BLB_DN[393] BLB_DN[394]
+ BLB_DN[395] BLB_DN[396] BLB_DN[397] BLB_DN[398] BLB_DN[399] BLB_DN[400]
+ BLB_DN[401] BLB_DN[402] BLB_DN[403] BLB_DN[404] BLB_DN[405] BLB_DN[406]
+ BLB_DN[407] BLB_DN[408] BLB_DN[409] BLB_DN[410] BLB_DN[411] BLB_DN[412]
+ BLB_DN[413] BLB_DN[414] BLB_DN[415] BLB_DN[416] BLB_DN[417] BLB_DN[418]
+ BLB_DN[419] BLB_DN[420] BLB_DN[421] BLB_DN[422] BLB_DN[423] BLB_DN[424]
+ BLB_DN[425] BLB_DN[426] BLB_DN[427] BLB_DN[428] BLB_DN[429] BLB_DN[430]
+ BLB_DN[431] BLB_DN[432] BLB_DN[433] BLB_DN[434] BLB_DN[435] BLB_DN[436]
+ BLB_DN[437] BLB_DN[438] BLB_DN[439] BLB_DN[440] BLB_DN[441] BLB_DN[442]
+ BLB_DN[443] BLB_DN[444] BLB_DN[445] BLB_DN[446] BLB_DN[447] BLB_DN[448]
+ BLB_DN[449] BLB_DN[450] BLB_DN[451] BLB_DN[452] BLB_DN[453] BLB_DN[454]
+ BLB_DN[455] BLB_DN[456] BLB_DN[457] BLB_DN[458] BLB_DN[459] BLB_DN[460]
+ BLB_DN[461] BLB_DN[462] BLB_DN[463] BLB_DN[464] BLB_DN[465] BLB_DN[466]
+ BLB_DN[467] BLB_DN[468] BLB_DN[469] BLB_DN[470] BLB_DN[471] BLB_DN[472]
+ BLB_DN[473] BLB_DN[474] BLB_DN[475] BLB_DN[476] BLB_DN[477] BLB_DN[478]
+ BLB_DN[479] BLB_DN[480] BLB_DN[481] BLB_DN[482] BLB_DN[483] BLB_DN[484]
+ BLB_DN[485] BLB_DN[486] BLB_DN[487] BLB_DN[488] BLB_DN[489] BLB_DN[490]
+ BLB_DN[491] BLB_DN[492] BLB_DN[493] BLB_DN[494] BLB_DN[495] BLB_DN[496]
+ BLB_DN[497] BLB_DN[498] BLB_DN[499] BLB_DN[500] BLB_DN[501] BLB_DN[502]
+ BLB_DN[503] BLB_DN[504] BLB_DN[505] BLB_DN[506] BLB_DN[507] BLB_DN[508]
+ BLB_DN[509] BLB_DN[510] BLB_DN[511] BLB_DN[512] BLB_DN[513] BLB_DN[514]
+ BLB_DN[515] BLB_DN[516] BLB_DN[517] BLB_DN[518] BLB_DN[519] BLB_DN[520]
+ BLB_DN[521] BLB_DN[522] BLB_DN[523] BLB_DN[524] BLB_DN[525] BLB_DN[526]
+ BLB_DN[527] BLB_DN[528] BLB_DN[529] BLB_DN[530] BLB_DN[531] BLB_DN[532]
+ BLB_DN[533] BLB_DN[534] BLB_DN[535] BLB_DN[536] BLB_DN[537] BLB_DN[538]
+ BLB_DN[539] BLB_DN[540] BLB_DN[541] BLB_DN[542] BLB_DN[543] BLB_DN[544]
+ BLB_DN[545] BLB_DN[546] BLB_DN[547] BLB_DN[548] BLB_DN[549] BLB_DN[550]
+ BLB_DN[551] BLB_DN[552] BLB_DN[553] BLB_DN[554] BLB_DN[555] BLB_DN[556]
+ BLB_DN[557] BLB_DN[558] BLB_DN[559] BLB_DN[560] BLB_DN[561] BLB_DN[562]
+ BLB_DN[563] BLB_DN[564] BLB_DN[565] BLB_DN[566] BLB_DN[567] BLB_DN[568]
+ BLB_DN[569] BLB_DN[570] BLB_DN[571] BLB_DN[572] BLB_DN[573] BLB_DN[574]
+ BLB_DN[575] BLB_UP[288] BLB_UP[289] BLB_UP[290] BLB_UP[291] BLB_UP[292]
+ BLB_UP[293] BLB_UP[294] BLB_UP[295] BLB_UP[296] BLB_UP[297] BLB_UP[298]
+ BLB_UP[299] BLB_UP[300] BLB_UP[301] BLB_UP[302] BLB_UP[303] BLB_UP[304]
+ BLB_UP[305] BLB_UP[306] BLB_UP[307] BLB_UP[308] BLB_UP[309] BLB_UP[310]
+ BLB_UP[311] BLB_UP[312] BLB_UP[313] BLB_UP[314] BLB_UP[315] BLB_UP[316]
+ BLB_UP[317] BLB_UP[318] BLB_UP[319] BLB_UP[320] BLB_UP[321] BLB_UP[322]
+ BLB_UP[323] BLB_UP[324] BLB_UP[325] BLB_UP[326] BLB_UP[327] BLB_UP[328]
+ BLB_UP[329] BLB_UP[330] BLB_UP[331] BLB_UP[332] BLB_UP[333] BLB_UP[334]
+ BLB_UP[335] BLB_UP[336] BLB_UP[337] BLB_UP[338] BLB_UP[339] BLB_UP[340]
+ BLB_UP[341] BLB_UP[342] BLB_UP[343] BLB_UP[344] BLB_UP[345] BLB_UP[346]
+ BLB_UP[347] BLB_UP[348] BLB_UP[349] BLB_UP[350] BLB_UP[351] BLB_UP[352]
+ BLB_UP[353] BLB_UP[354] BLB_UP[355] BLB_UP[356] BLB_UP[357] BLB_UP[358]
+ BLB_UP[359] BLB_UP[360] BLB_UP[361] BLB_UP[362] BLB_UP[363] BLB_UP[364]
+ BLB_UP[365] BLB_UP[366] BLB_UP[367] BLB_UP[368] BLB_UP[369] BLB_UP[370]
+ BLB_UP[371] BLB_UP[372] BLB_UP[373] BLB_UP[374] BLB_UP[375] BLB_UP[376]
+ BLB_UP[377] BLB_UP[378] BLB_UP[379] BLB_UP[380] BLB_UP[381] BLB_UP[382]
+ BLB_UP[383] BLB_UP[384] BLB_UP[385] BLB_UP[386] BLB_UP[387] BLB_UP[388]
+ BLB_UP[389] BLB_UP[390] BLB_UP[391] BLB_UP[392] BLB_UP[393] BLB_UP[394]
+ BLB_UP[395] BLB_UP[396] BLB_UP[397] BLB_UP[398] BLB_UP[399] BLB_UP[400]
+ BLB_UP[401] BLB_UP[402] BLB_UP[403] BLB_UP[404] BLB_UP[405] BLB_UP[406]
+ BLB_UP[407] BLB_UP[408] BLB_UP[409] BLB_UP[410] BLB_UP[411] BLB_UP[412]
+ BLB_UP[413] BLB_UP[414] BLB_UP[415] BLB_UP[416] BLB_UP[417] BLB_UP[418]
+ BLB_UP[419] BLB_UP[420] BLB_UP[421] BLB_UP[422] BLB_UP[423] BLB_UP[424]
+ BLB_UP[425] BLB_UP[426] BLB_UP[427] BLB_UP[428] BLB_UP[429] BLB_UP[430]
+ BLB_UP[431] BLB_UP[432] BLB_UP[433] BLB_UP[434] BLB_UP[435] BLB_UP[436]
+ BLB_UP[437] BLB_UP[438] BLB_UP[439] BLB_UP[440] BLB_UP[441] BLB_UP[442]
+ BLB_UP[443] BLB_UP[444] BLB_UP[445] BLB_UP[446] BLB_UP[447] BLB_UP[448]
+ BLB_UP[449] BLB_UP[450] BLB_UP[451] BLB_UP[452] BLB_UP[453] BLB_UP[454]
+ BLB_UP[455] BLB_UP[456] BLB_UP[457] BLB_UP[458] BLB_UP[459] BLB_UP[460]
+ BLB_UP[461] BLB_UP[462] BLB_UP[463] BLB_UP[464] BLB_UP[465] BLB_UP[466]
+ BLB_UP[467] BLB_UP[468] BLB_UP[469] BLB_UP[470] BLB_UP[471] BLB_UP[472]
+ BLB_UP[473] BLB_UP[474] BLB_UP[475] BLB_UP[476] BLB_UP[477] BLB_UP[478]
+ BLB_UP[479] BLB_UP[480] BLB_UP[481] BLB_UP[482] BLB_UP[483] BLB_UP[484]
+ BLB_UP[485] BLB_UP[486] BLB_UP[487] BLB_UP[488] BLB_UP[489] BLB_UP[490]
+ BLB_UP[491] BLB_UP[492] BLB_UP[493] BLB_UP[494] BLB_UP[495] BLB_UP[496]
+ BLB_UP[497] BLB_UP[498] BLB_UP[499] BLB_UP[500] BLB_UP[501] BLB_UP[502]
+ BLB_UP[503] BLB_UP[504] BLB_UP[505] BLB_UP[506] BLB_UP[507] BLB_UP[508]
+ BLB_UP[509] BLB_UP[510] BLB_UP[511] BLB_UP[512] BLB_UP[513] BLB_UP[514]
+ BLB_UP[515] BLB_UP[516] BLB_UP[517] BLB_UP[518] BLB_UP[519] BLB_UP[520]
+ BLB_UP[521] BLB_UP[522] BLB_UP[523] BLB_UP[524] BLB_UP[525] BLB_UP[526]
+ BLB_UP[527] BLB_UP[528] BLB_UP[529] BLB_UP[530] BLB_UP[531] BLB_UP[532]
+ BLB_UP[533] BLB_UP[534] BLB_UP[535] BLB_UP[536] BLB_UP[537] BLB_UP[538]
+ BLB_UP[539] BLB_UP[540] BLB_UP[541] BLB_UP[542] BLB_UP[543] BLB_UP[544]
+ BLB_UP[545] BLB_UP[546] BLB_UP[547] BLB_UP[548] BLB_UP[549] BLB_UP[550]
+ BLB_UP[551] BLB_UP[552] BLB_UP[553] BLB_UP[554] BLB_UP[555] BLB_UP[556]
+ BLB_UP[557] BLB_UP[558] BLB_UP[559] BLB_UP[560] BLB_UP[561] BLB_UP[562]
+ BLB_UP[563] BLB_UP[564] BLB_UP[565] BLB_UP[566] BLB_UP[567] BLB_UP[568]
+ BLB_UP[569] BLB_UP[570] BLB_UP[571] BLB_UP[572] BLB_UP[573] BLB_UP[574]
+ BLB_UP[575] BLEQ_DN BLEQ_UP BL_DN[288] BL_DN[289] BL_DN[290] BL_DN[291]
+ BL_DN[292] BL_DN[293] BL_DN[294] BL_DN[295] BL_DN[296] BL_DN[297] BL_DN[298]
+ BL_DN[299] BL_DN[300] BL_DN[301] BL_DN[302] BL_DN[303] BL_DN[304] BL_DN[305]
+ BL_DN[306] BL_DN[307] BL_DN[308] BL_DN[309] BL_DN[310] BL_DN[311] BL_DN[312]
+ BL_DN[313] BL_DN[314] BL_DN[315] BL_DN[316] BL_DN[317] BL_DN[318] BL_DN[319]
+ BL_DN[320] BL_DN[321] BL_DN[322] BL_DN[323] BL_DN[324] BL_DN[325] BL_DN[326]
+ BL_DN[327] BL_DN[328] BL_DN[329] BL_DN[330] BL_DN[331] BL_DN[332] BL_DN[333]
+ BL_DN[334] BL_DN[335] BL_DN[336] BL_DN[337] BL_DN[338] BL_DN[339] BL_DN[340]
+ BL_DN[341] BL_DN[342] BL_DN[343] BL_DN[344] BL_DN[345] BL_DN[346] BL_DN[347]
+ BL_DN[348] BL_DN[349] BL_DN[350] BL_DN[351] BL_DN[352] BL_DN[353] BL_DN[354]
+ BL_DN[355] BL_DN[356] BL_DN[357] BL_DN[358] BL_DN[359] BL_DN[360] BL_DN[361]
+ BL_DN[362] BL_DN[363] BL_DN[364] BL_DN[365] BL_DN[366] BL_DN[367] BL_DN[368]
+ BL_DN[369] BL_DN[370] BL_DN[371] BL_DN[372] BL_DN[373] BL_DN[374] BL_DN[375]
+ BL_DN[376] BL_DN[377] BL_DN[378] BL_DN[379] BL_DN[380] BL_DN[381] BL_DN[382]
+ BL_DN[383] BL_DN[384] BL_DN[385] BL_DN[386] BL_DN[387] BL_DN[388] BL_DN[389]
+ BL_DN[390] BL_DN[391] BL_DN[392] BL_DN[393] BL_DN[394] BL_DN[395] BL_DN[396]
+ BL_DN[397] BL_DN[398] BL_DN[399] BL_DN[400] BL_DN[401] BL_DN[402] BL_DN[403]
+ BL_DN[404] BL_DN[405] BL_DN[406] BL_DN[407] BL_DN[408] BL_DN[409] BL_DN[410]
+ BL_DN[411] BL_DN[412] BL_DN[413] BL_DN[414] BL_DN[415] BL_DN[416] BL_DN[417]
+ BL_DN[418] BL_DN[419] BL_DN[420] BL_DN[421] BL_DN[422] BL_DN[423] BL_DN[424]
+ BL_DN[425] BL_DN[426] BL_DN[427] BL_DN[428] BL_DN[429] BL_DN[430] BL_DN[431]
+ BL_DN[432] BL_DN[433] BL_DN[434] BL_DN[435] BL_DN[436] BL_DN[437] BL_DN[438]
+ BL_DN[439] BL_DN[440] BL_DN[441] BL_DN[442] BL_DN[443] BL_DN[444] BL_DN[445]
+ BL_DN[446] BL_DN[447] BL_DN[448] BL_DN[449] BL_DN[450] BL_DN[451] BL_DN[452]
+ BL_DN[453] BL_DN[454] BL_DN[455] BL_DN[456] BL_DN[457] BL_DN[458] BL_DN[459]
+ BL_DN[460] BL_DN[461] BL_DN[462] BL_DN[463] BL_DN[464] BL_DN[465] BL_DN[466]
+ BL_DN[467] BL_DN[468] BL_DN[469] BL_DN[470] BL_DN[471] BL_DN[472] BL_DN[473]
+ BL_DN[474] BL_DN[475] BL_DN[476] BL_DN[477] BL_DN[478] BL_DN[479] BL_DN[480]
+ BL_DN[481] BL_DN[482] BL_DN[483] BL_DN[484] BL_DN[485] BL_DN[486] BL_DN[487]
+ BL_DN[488] BL_DN[489] BL_DN[490] BL_DN[491] BL_DN[492] BL_DN[493] BL_DN[494]
+ BL_DN[495] BL_DN[496] BL_DN[497] BL_DN[498] BL_DN[499] BL_DN[500] BL_DN[501]
+ BL_DN[502] BL_DN[503] BL_DN[504] BL_DN[505] BL_DN[506] BL_DN[507] BL_DN[508]
+ BL_DN[509] BL_DN[510] BL_DN[511] BL_DN[512] BL_DN[513] BL_DN[514] BL_DN[515]
+ BL_DN[516] BL_DN[517] BL_DN[518] BL_DN[519] BL_DN[520] BL_DN[521] BL_DN[522]
+ BL_DN[523] BL_DN[524] BL_DN[525] BL_DN[526] BL_DN[527] BL_DN[528] BL_DN[529]
+ BL_DN[530] BL_DN[531] BL_DN[532] BL_DN[533] BL_DN[534] BL_DN[535] BL_DN[536]
+ BL_DN[537] BL_DN[538] BL_DN[539] BL_DN[540] BL_DN[541] BL_DN[542] BL_DN[543]
+ BL_DN[544] BL_DN[545] BL_DN[546] BL_DN[547] BL_DN[548] BL_DN[549] BL_DN[550]
+ BL_DN[551] BL_DN[552] BL_DN[553] BL_DN[554] BL_DN[555] BL_DN[556] BL_DN[557]
+ BL_DN[558] BL_DN[559] BL_DN[560] BL_DN[561] BL_DN[562] BL_DN[563] BL_DN[564]
+ BL_DN[565] BL_DN[566] BL_DN[567] BL_DN[568] BL_DN[569] BL_DN[570] BL_DN[571]
+ BL_DN[572] BL_DN[573] BL_DN[574] BL_DN[575] BL_UP[288] BL_UP[289] BL_UP[290]
+ BL_UP[291] BL_UP[292] BL_UP[293] BL_UP[294] BL_UP[295] BL_UP[296] BL_UP[297]
+ BL_UP[298] BL_UP[299] BL_UP[300] BL_UP[301] BL_UP[302] BL_UP[303] BL_UP[304]
+ BL_UP[305] BL_UP[306] BL_UP[307] BL_UP[308] BL_UP[309] BL_UP[310] BL_UP[311]
+ BL_UP[312] BL_UP[313] BL_UP[314] BL_UP[315] BL_UP[316] BL_UP[317] BL_UP[318]
+ BL_UP[319] BL_UP[320] BL_UP[321] BL_UP[322] BL_UP[323] BL_UP[324] BL_UP[325]
+ BL_UP[326] BL_UP[327] BL_UP[328] BL_UP[329] BL_UP[330] BL_UP[331] BL_UP[332]
+ BL_UP[333] BL_UP[334] BL_UP[335] BL_UP[336] BL_UP[337] BL_UP[338] BL_UP[339]
+ BL_UP[340] BL_UP[341] BL_UP[342] BL_UP[343] BL_UP[344] BL_UP[345] BL_UP[346]
+ BL_UP[347] BL_UP[348] BL_UP[349] BL_UP[350] BL_UP[351] BL_UP[352] BL_UP[353]
+ BL_UP[354] BL_UP[355] BL_UP[356] BL_UP[357] BL_UP[358] BL_UP[359] BL_UP[360]
+ BL_UP[361] BL_UP[362] BL_UP[363] BL_UP[364] BL_UP[365] BL_UP[366] BL_UP[367]
+ BL_UP[368] BL_UP[369] BL_UP[370] BL_UP[371] BL_UP[372] BL_UP[373] BL_UP[374]
+ BL_UP[375] BL_UP[376] BL_UP[377] BL_UP[378] BL_UP[379] BL_UP[380] BL_UP[381]
+ BL_UP[382] BL_UP[383] BL_UP[384] BL_UP[385] BL_UP[386] BL_UP[387] BL_UP[388]
+ BL_UP[389] BL_UP[390] BL_UP[391] BL_UP[392] BL_UP[393] BL_UP[394] BL_UP[395]
+ BL_UP[396] BL_UP[397] BL_UP[398] BL_UP[399] BL_UP[400] BL_UP[401] BL_UP[402]
+ BL_UP[403] BL_UP[404] BL_UP[405] BL_UP[406] BL_UP[407] BL_UP[408] BL_UP[409]
+ BL_UP[410] BL_UP[411] BL_UP[412] BL_UP[413] BL_UP[414] BL_UP[415] BL_UP[416]
+ BL_UP[417] BL_UP[418] BL_UP[419] BL_UP[420] BL_UP[421] BL_UP[422] BL_UP[423]
+ BL_UP[424] BL_UP[425] BL_UP[426] BL_UP[427] BL_UP[428] BL_UP[429] BL_UP[430]
+ BL_UP[431] BL_UP[432] BL_UP[433] BL_UP[434] BL_UP[435] BL_UP[436] BL_UP[437]
+ BL_UP[438] BL_UP[439] BL_UP[440] BL_UP[441] BL_UP[442] BL_UP[443] BL_UP[444]
+ BL_UP[445] BL_UP[446] BL_UP[447] BL_UP[448] BL_UP[449] BL_UP[450] BL_UP[451]
+ BL_UP[452] BL_UP[453] BL_UP[454] BL_UP[455] BL_UP[456] BL_UP[457] BL_UP[458]
+ BL_UP[459] BL_UP[460] BL_UP[461] BL_UP[462] BL_UP[463] BL_UP[464] BL_UP[465]
+ BL_UP[466] BL_UP[467] BL_UP[468] BL_UP[469] BL_UP[470] BL_UP[471] BL_UP[472]
+ BL_UP[473] BL_UP[474] BL_UP[475] BL_UP[476] BL_UP[477] BL_UP[478] BL_UP[479]
+ BL_UP[480] BL_UP[481] BL_UP[482] BL_UP[483] BL_UP[484] BL_UP[485] BL_UP[486]
+ BL_UP[487] BL_UP[488] BL_UP[489] BL_UP[490] BL_UP[491] BL_UP[492] BL_UP[493]
+ BL_UP[494] BL_UP[495] BL_UP[496] BL_UP[497] BL_UP[498] BL_UP[499] BL_UP[500]
+ BL_UP[501] BL_UP[502] BL_UP[503] BL_UP[504] BL_UP[505] BL_UP[506] BL_UP[507]
+ BL_UP[508] BL_UP[509] BL_UP[510] BL_UP[511] BL_UP[512] BL_UP[513] BL_UP[514]
+ BL_UP[515] BL_UP[516] BL_UP[517] BL_UP[518] BL_UP[519] BL_UP[520] BL_UP[521]
+ BL_UP[522] BL_UP[523] BL_UP[524] BL_UP[525] BL_UP[526] BL_UP[527] BL_UP[528]
+ BL_UP[529] BL_UP[530] BL_UP[531] BL_UP[532] BL_UP[533] BL_UP[534] BL_UP[535]
+ BL_UP[536] BL_UP[537] BL_UP[538] BL_UP[539] BL_UP[540] BL_UP[541] BL_UP[542]
+ BL_UP[543] BL_UP[544] BL_UP[545] BL_UP[546] BL_UP[547] BL_UP[548] BL_UP[549]
+ BL_UP[550] BL_UP[551] BL_UP[552] BL_UP[553] BL_UP[554] BL_UP[555] BL_UP[556]
+ BL_UP[557] BL_UP[558] BL_UP[559] BL_UP[560] BL_UP[561] BL_UP[562] BL_UP[563]
+ BL_UP[564] BL_UP[565] BL_UP[566] BL_UP[567] BL_UP[568] BL_UP[569] BL_UP[570]
+ BL_UP[571] BL_UP[572] BL_UP[573] BL_UP[574] BL_UP[575] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[18] GBLB[19] GBLB[20]
+ GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28]
+ GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[18] GW[19]
+ GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30]
+ GW[31] GW[32] GW[33] GW[34] GW[35] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22]
+ GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31]
+ GWB[32] GWB[33] GWB[34] GWB[35] LIOPD LIOPD PDOXR RE SAEB VXDDAI VDDI VSSI WE
+ YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6]
+ Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ S1BSVTSWSO8000Y24_LIO_R_SD
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_BANK_F_UP_REP GBL[0] GBL[1] GBL[2] GBL[3] GBL[4]
+ GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14]
+ GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23]
+ GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32]
+ GBL[33] GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5]
+ GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14]
+ GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22]
+ GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30]
+ GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2]
+ GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12]
+ GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21]
+ GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30]
+ GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] DSLP_BUF SLP_LCTRL SLP_LCTRL_REP RE WE
+ VXDDHD WLP_SAE DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1[0] DEC_X1[1]
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] YL[1]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] VXDDAI VDDI VSSI WLP_SAE_TK TK
XLIO_MCB_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] VXDDAI LIOPD WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7]
+ WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18]
+ WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29]
+ WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40]
+ WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51]
+ WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62]
+ WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73]
+ WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84]
+ WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95]
+ WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105]
+ WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114]
+ WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123]
+ WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] WL[132]
+ WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141]
+ WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150]
+ WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159]
+ WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168]
+ WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177]
+ WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186]
+ WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] WL[195]
+ WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204]
+ WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213]
+ WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222]
+ WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231]
+ WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240]
+ WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249]
+ WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] WL[258]
+ WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] WL[267]
+ WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] WL[276]
+ WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] WL[285]
+ WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] WL[294]
+ WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] WL[303]
+ WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] WL[312]
+ WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] WL[321]
+ WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] WL[330]
+ WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] WL[339]
+ WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] WL[348]
+ WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] WL[357]
+ WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] WL[366]
+ WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] WL[375]
+ WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] WL[383] WL[384]
+ WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] WL[392] WL[393]
+ WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] WL[401] WL[402]
+ WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] WL[410] WL[411]
+ WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] WL[419] WL[420]
+ WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] WL[428] WL[429]
+ WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] WL[437] WL[438]
+ WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] WL[446] WL[447]
+ WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] WL[455] WL[456]
+ WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] WL[464] WL[465]
+ WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] WL[473] WL[474]
+ WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] WL[482] WL[483]
+ WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] WL[491] WL[492]
+ WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] WL[500] WL[501]
+ WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] WL[509] WL[510]
+ WL[511] BLEQ_DN BLEQ_UP GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8]
+ GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19]
+ GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30]
+ GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5]
+ GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15]
+ GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24]
+ GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33]
+ GWB[34] GWB[35] RE_LIO SAEB WE_LIO DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2]
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0]
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6]
+ DEC_Y_UP[7] YL_LIO[0] YL_LIO[1] VDDI VSSI S1BSVTSWSO8000Y24_LIO_MCB_F
XLCTRL_S_M16_SD BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1]
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4]
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4]
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3]
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1]
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7]
+ DSLP_BUF LIOPD RE RE_LIO SAEB SLP_LCTRL TK VXDDHD VDDI VSSI WE WE_LIO
+ WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2]
+ WLPY_UP[3] WLP_SAE WLP_SAE_TK YL[0] YL[1] YL_LIO[0] YL_LIO[1]
+ S1BSVTSWSO8000Y24_LCTRL_S_M16_SD
XXDRV_STRAPD0 VXDDHD VDDI VSSI WLPY_DN[0] WLPY_DNB[0]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_SHA_0 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD0 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[0] WL[1]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_1 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD0 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[2] WL[3]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS1 DEC_X1[0] SH_NPD0 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_2 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD1 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[4] WL[5]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_3 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD1 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[6] WL[7]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS3 DEC_X1[0] SH_NPD1 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_4 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD2 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[8] WL[9]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_5 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD2 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[10] WL[11]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS5 DEC_X1[1] SH_NPD2 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_6 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD3 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[12] WL[13]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_7 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD3 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[14] WL[15]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS7 DEC_X1[1] SH_NPD3 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_8 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD4 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[16] WL[17]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_9 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD4 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[18] WL[19]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS9 DEC_X1[2] SH_NPD4 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_10 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD5 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[20] WL[21]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_11 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD5 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[22] WL[23]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS11 DEC_X1[2] SH_NPD5 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_12 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD6 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[24] WL[25]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_13 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD6 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[26] WL[27]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS13 DEC_X1[3] SH_NPD6 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_14 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD7 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[28] WL[29]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_15 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD7 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[30] WL[31]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS15 DEC_X1[3] SH_NPD7 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_16 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD8 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[32] WL[33]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_17 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD8 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[34] WL[35]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS17 DEC_X1[4] SH_NPD8 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_18 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD9 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[36] WL[37]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_19 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD9 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[38] WL[39]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS19 DEC_X1[4] SH_NPD9 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_20 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD10 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[40] WL[41]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_21 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD10 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[42] WL[43]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS21 DEC_X1[5] SH_NPD10 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_22 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD11 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[44] WL[45]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_23 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD11 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[46] WL[47]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS23 DEC_X1[5] SH_NPD11 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_24 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD12 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[48] WL[49]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_25 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD12 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[50] WL[51]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS25 DEC_X1[6] SH_NPD12 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_26 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD13 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[52] WL[53]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_27 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD13 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[54] WL[55]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS27 DEC_X1[6] SH_NPD13 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_28 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD14 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[56] WL[57]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_29 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD14 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[58] WL[59]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS29 DEC_X1[7] SH_NPD14 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_30 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD15 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[60] WL[61]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_31 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD15 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[62] WL[63]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS31 DEC_X1[7] SH_NPD15 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPD1 VXDDHD VDDI VSSI WLPY_DN[1] WLPY_DNB[1]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_SHA_32 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD16 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[64] WL[65]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_33 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD16 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[66] WL[67]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS33 DEC_X1[0] SH_NPD16 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_34 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD17 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[68] WL[69]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_35 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD17 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[70] WL[71]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS35 DEC_X1[0] SH_NPD17 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_36 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD18 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[72] WL[73]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_37 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD18 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[74] WL[75]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS37 DEC_X1[1] SH_NPD18 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_38 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD19 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[76] WL[77]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_39 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD19 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[78] WL[79]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS39 DEC_X1[1] SH_NPD19 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_40 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD20 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[80] WL[81]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_41 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD20 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[82] WL[83]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS41 DEC_X1[2] SH_NPD20 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_42 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD21 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[84] WL[85]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_43 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD21 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[86] WL[87]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS43 DEC_X1[2] SH_NPD21 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_44 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD22 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[88] WL[89]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_45 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD22 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[90] WL[91]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS45 DEC_X1[3] SH_NPD22 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_46 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD23 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[92] WL[93]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_47 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD23 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[94] WL[95]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS47 DEC_X1[3] SH_NPD23 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_48 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD24 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[96] WL[97]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_49 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD24 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[98] WL[99]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS49 DEC_X1[4] SH_NPD24 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_50 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD25 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[100] WL[101]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_51 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD25 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[102] WL[103]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS51 DEC_X1[4] SH_NPD25 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_52 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD26 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[104] WL[105]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_53 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD26 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[106] WL[107]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS53 DEC_X1[5] SH_NPD26 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_54 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD27 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[108] WL[109]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_55 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD27 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[110] WL[111]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS55 DEC_X1[5] SH_NPD27 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_56 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD28 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[112] WL[113]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_57 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD28 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[114] WL[115]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS57 DEC_X1[6] SH_NPD28 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_58 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD29 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[116] WL[117]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_59 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD29 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[118] WL[119]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS59 DEC_X1[6] SH_NPD29 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_60 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD30 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[120] WL[121]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_61 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD30 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[122] WL[123]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS61 DEC_X1[7] SH_NPD30 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_62 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD31 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[124] WL[125]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_63 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD31 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[126] WL[127]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS63 DEC_X1[7] SH_NPD31 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPD2 VXDDHD VDDI VSSI WLPY_DN[2] WLPY_DNB[2]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_SHA_64 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD32 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[128] WL[129]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_65 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD32 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[130] WL[131]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS65 DEC_X1[0] SH_NPD32 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_66 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD33 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[132] WL[133]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_67 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD33 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[134] WL[135]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS67 DEC_X1[0] SH_NPD33 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_68 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD34 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[136] WL[137]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_69 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD34 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[138] WL[139]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS69 DEC_X1[1] SH_NPD34 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_70 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD35 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[140] WL[141]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_71 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD35 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[142] WL[143]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS71 DEC_X1[1] SH_NPD35 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_72 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD36 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[144] WL[145]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_73 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD36 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[146] WL[147]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS73 DEC_X1[2] SH_NPD36 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_74 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD37 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[148] WL[149]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_75 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD37 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[150] WL[151]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS75 DEC_X1[2] SH_NPD37 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_76 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD38 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[152] WL[153]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_77 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD38 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[154] WL[155]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS77 DEC_X1[3] SH_NPD38 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_78 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD39 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[156] WL[157]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_79 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD39 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[158] WL[159]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS79 DEC_X1[3] SH_NPD39 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_80 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD40 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[160] WL[161]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_81 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD40 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[162] WL[163]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS81 DEC_X1[4] SH_NPD40 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_82 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD41 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[164] WL[165]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_83 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD41 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[166] WL[167]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS83 DEC_X1[4] SH_NPD41 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_84 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD42 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[168] WL[169]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_85 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD42 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[170] WL[171]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS85 DEC_X1[5] SH_NPD42 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_86 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD43 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[172] WL[173]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_87 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD43 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[174] WL[175]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS87 DEC_X1[5] SH_NPD43 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_88 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD44 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[176] WL[177]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_89 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD44 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[178] WL[179]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS89 DEC_X1[6] SH_NPD44 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_90 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD45 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[180] WL[181]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_91 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD45 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[182] WL[183]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS91 DEC_X1[6] SH_NPD45 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_92 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD46 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[184] WL[185]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_93 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD46 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[186] WL[187]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS93 DEC_X1[7] SH_NPD46 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_94 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD47 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[188] WL[189]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_95 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD47 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[190] WL[191]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS95 DEC_X1[7] SH_NPD47 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPD3 VXDDHD VDDI VSSI WLPY_DN[3] WLPY_DNB[3]
+ S1BSVTSWSO8000Y24_XDRV_STRAP_LCNT
XXDRV_LA512_SHA_96 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD48 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[192] WL[193]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_97 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD48 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[194] WL[195]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS97 DEC_X1[0] SH_NPD48 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_98 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD49 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[196] WL[197]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_99 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD49 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[198] WL[199]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS99 DEC_X1[0] SH_NPD49 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_100 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD50 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[200] WL[201]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_101 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD50 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[202] WL[203]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS101 DEC_X1[1] SH_NPD50 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_102 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD51 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[204] WL[205]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_103 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD51 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[206] WL[207]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS103 DEC_X1[1] SH_NPD51 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_104 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD52 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[208] WL[209]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_105 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD52 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[210] WL[211]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS105 DEC_X1[2] SH_NPD52 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_106 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD53 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[212] WL[213]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_107 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD53 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[214] WL[215]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS107 DEC_X1[2] SH_NPD53 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_108 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD54 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[216] WL[217]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_109 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD54 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[218] WL[219]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS109 DEC_X1[3] SH_NPD54 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_110 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD55 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[220] WL[221]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_111 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD55 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[222] WL[223]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS111 DEC_X1[3] SH_NPD55 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_112 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD56 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[224] WL[225]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_113 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD56 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[226] WL[227]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS113 DEC_X1[4] SH_NPD56 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_114 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD57 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[228] WL[229]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_115 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD57 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[230] WL[231]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS115 DEC_X1[4] SH_NPD57 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_116 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD58 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[232] WL[233]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_117 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD58 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[234] WL[235]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS117 DEC_X1[5] SH_NPD58 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_118 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD59 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[236] WL[237]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_119 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD59 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[238] WL[239]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS119 DEC_X1[5] SH_NPD59 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_120 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD60 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[240] WL[241]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_121 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD60 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[242] WL[243]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS121 DEC_X1[6] SH_NPD60 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_122 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD61 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[244] WL[245]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_123 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD61 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[246] WL[247]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS123 DEC_X1[6] SH_NPD61 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_124 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD62 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[248] WL[249]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_125 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD62 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[250] WL[251]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS125 DEC_X1[7] SH_NPD62 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_126 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD63 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[252] WL[253]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_127 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD63 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[254] WL[255]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS127 DEC_X1[7] SH_NPD63 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPU0 VXDDHD VDDI VSSI WLPY_UP[0] WLPY_UPB[0]
+ S1BSVTSWSO8000Y24_XDRV_STRAP_LCNT
XXDRV_LA512_NOR_SHA_128 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD64 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[256] WL[257] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_129 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD64 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[258] WL[259] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS129 DEC_X1_REP[0] SH_NPD64 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_130 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD65 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[260] WL[261] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_131 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD65 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[262] WL[263] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS131 DEC_X1_REP[0] SH_NPD65 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_132 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD66 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[264] WL[265] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_133 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD66 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[266] WL[267] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS133 DEC_X1_REP[1] SH_NPD66 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_134 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD67 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[268] WL[269] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_135 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD67 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[270] WL[271] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS135 DEC_X1_REP[1] SH_NPD67 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_136 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD68 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[272] WL[273] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_137 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD68 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[274] WL[275] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS137 DEC_X1_REP[2] SH_NPD68 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_138 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD69 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[276] WL[277] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_139 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD69 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[278] WL[279] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS139 DEC_X1_REP[2] SH_NPD69 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_140 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD70 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[280] WL[281] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_141 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD70 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[282] WL[283] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS141 DEC_X1_REP[3] SH_NPD70 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_142 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD71 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[284] WL[285] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_143 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD71 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[286] WL[287] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS143 DEC_X1_REP[3] SH_NPD71 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_144 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD72 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[288] WL[289] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_145 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD72 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[290] WL[291] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS145 DEC_X1_REP[4] SH_NPD72 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_146 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD73 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[292] WL[293] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_147 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD73 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[294] WL[295] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS147 DEC_X1_REP[4] SH_NPD73 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_148 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD74 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[296] WL[297] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_149 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD74 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[298] WL[299] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS149 DEC_X1_REP[5] SH_NPD74 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_150 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD75 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[300] WL[301] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_151 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD75 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[302] WL[303] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS151 DEC_X1_REP[5] SH_NPD75 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_152 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD76 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[304] WL[305] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_153 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD76 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[306] WL[307] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS153 DEC_X1_REP[6] SH_NPD76 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_154 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD77 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[308] WL[309] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_155 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD77 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[310] WL[311] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS155 DEC_X1_REP[6] SH_NPD77 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_156 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD78 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[312] WL[313] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_157 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD78 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[314] WL[315] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS157 DEC_X1_REP[7] SH_NPD78 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_158 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD79 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[316] WL[317] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_159 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD79 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[318] WL[319] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS159 DEC_X1_REP[7] SH_NPD79 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_STRAPU1 VXDDHD VDDI VSSI WLPY_UP[1] WLPY_UPB[1]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_NOR_SHA_160 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD80 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[320] WL[321] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_161 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD80 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[322] WL[323] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS161 DEC_X1_REP[0] SH_NPD80 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_162 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD81 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[324] WL[325] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_163 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD81 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[326] WL[327] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS163 DEC_X1_REP[0] SH_NPD81 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_164 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD82 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[328] WL[329] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_165 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD82 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[330] WL[331] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS165 DEC_X1_REP[1] SH_NPD82 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_166 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD83 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[332] WL[333] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_167 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD83 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[334] WL[335] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS167 DEC_X1_REP[1] SH_NPD83 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_168 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD84 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[336] WL[337] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_169 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD84 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[338] WL[339] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS169 DEC_X1_REP[2] SH_NPD84 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_170 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD85 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[340] WL[341] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_171 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD85 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[342] WL[343] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS171 DEC_X1_REP[2] SH_NPD85 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_172 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD86 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[344] WL[345] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_173 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD86 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[346] WL[347] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS173 DEC_X1_REP[3] SH_NPD86 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_174 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD87 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[348] WL[349] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_175 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD87 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[350] WL[351] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS175 DEC_X1_REP[3] SH_NPD87 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_176 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD88 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[352] WL[353] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_177 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD88 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[354] WL[355] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS177 DEC_X1_REP[4] SH_NPD88 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_178 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD89 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[356] WL[357] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_179 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD89 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[358] WL[359] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS179 DEC_X1_REP[4] SH_NPD89 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_180 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD90 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[360] WL[361] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_181 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD90 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[362] WL[363] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS181 DEC_X1_REP[5] SH_NPD90 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_182 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD91 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[364] WL[365] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_183 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD91 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[366] WL[367] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS183 DEC_X1_REP[5] SH_NPD91 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_184 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD92 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[368] WL[369] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_185 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD92 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[370] WL[371] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS185 DEC_X1_REP[6] SH_NPD92 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_186 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD93 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[372] WL[373] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_187 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD93 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[374] WL[375] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS187 DEC_X1_REP[6] SH_NPD93 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_188 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD94 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[376] WL[377] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_189 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD94 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[378] WL[379] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS189 DEC_X1_REP[7] SH_NPD94 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_190 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD95 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[380] WL[381] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_191 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD95 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[382] WL[383] WLPY_UP[1]
+ WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS191 DEC_X1_REP[7] SH_NPD95 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_STRAPU2 VXDDHD VDDI VSSI WLPY_UP[2] WLPY_UPB[2]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_NOR_SHA_192 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD96 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[384] WL[385] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_193 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD96 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[386] WL[387] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS193 DEC_X1_REP[0] SH_NPD96 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_194 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD97 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[388] WL[389] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_195 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD97 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[390] WL[391] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS195 DEC_X1_REP[0] SH_NPD97 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_196 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD98 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[392] WL[393] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_197 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD98 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[394] WL[395] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS197 DEC_X1_REP[1] SH_NPD98 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_198 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD99 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[396] WL[397] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_199 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD99 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[398] WL[399] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS199 DEC_X1_REP[1] SH_NPD99 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_200 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD100 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[400] WL[401] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_201 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD100 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[402] WL[403] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS201 DEC_X1_REP[2] SH_NPD100 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_202 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD101 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[404] WL[405] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_203 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD101 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[406] WL[407] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS203 DEC_X1_REP[2] SH_NPD101 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_204 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD102 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[408] WL[409] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_205 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD102 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[410] WL[411] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS205 DEC_X1_REP[3] SH_NPD102 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_206 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD103 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[412] WL[413] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_207 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD103 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[414] WL[415] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS207 DEC_X1_REP[3] SH_NPD103 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_208 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD104 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[416] WL[417] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_209 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD104 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[418] WL[419] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS209 DEC_X1_REP[4] SH_NPD104 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_210 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD105 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[420] WL[421] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_211 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD105 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[422] WL[423] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS211 DEC_X1_REP[4] SH_NPD105 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_212 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD106 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[424] WL[425] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_213 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD106 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[426] WL[427] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS213 DEC_X1_REP[5] SH_NPD106 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_214 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD107 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[428] WL[429] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_215 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD107 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[430] WL[431] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS215 DEC_X1_REP[5] SH_NPD107 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_216 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD108 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[432] WL[433] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_217 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD108 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[434] WL[435] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS217 DEC_X1_REP[6] SH_NPD108 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_218 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD109 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[436] WL[437] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_219 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD109 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[438] WL[439] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS219 DEC_X1_REP[6] SH_NPD109 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_220 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD110 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[440] WL[441] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_221 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD110 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[442] WL[443] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS221 DEC_X1_REP[7] SH_NPD110 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_222 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD111 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[444] WL[445] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_223 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD111 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[446] WL[447] WLPY_UP[2]
+ WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS223 DEC_X1_REP[7] SH_NPD111 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_STRAPU3 VXDDHD VDDI VSSI WLPY_UP[3] WLPY_UPB[3]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_NOR_SHA_224 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD112 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[448] WL[449] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_225 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD112 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[450] WL[451] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS225 DEC_X1_REP[0] SH_NPD112 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_226 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD113 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[452] WL[453] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_227 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD113 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[454] WL[455] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS227 DEC_X1_REP[0] SH_NPD113 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_228 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD114 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[456] WL[457] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_229 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD114 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[458] WL[459] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS229 DEC_X1_REP[1] SH_NPD114 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_230 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD115 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[460] WL[461] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_231 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[1]
+ DEC_X1_REP[0] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD115 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[462] WL[463] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS231 DEC_X1_REP[1] SH_NPD115 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_232 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD116 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[464] WL[465] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_233 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD116 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[466] WL[467] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS233 DEC_X1_REP[2] SH_NPD116 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_234 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD117 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[468] WL[469] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_235 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[2]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD117 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[470] WL[471] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS235 DEC_X1_REP[2] SH_NPD117 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_236 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD118 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[472] WL[473] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_237 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD118 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[474] WL[475] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS237 DEC_X1_REP[3] SH_NPD118 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_238 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD119 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[476] WL[477] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_239 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[3]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD119 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[478] WL[479] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS239 DEC_X1_REP[3] SH_NPD119 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_240 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD120 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[480] WL[481] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_241 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD120 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[482] WL[483] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS241 DEC_X1_REP[4] SH_NPD120 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_242 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD121 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[484] WL[485] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_243 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[4]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD121 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[486] WL[487] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS243 DEC_X1_REP[4] SH_NPD121 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_244 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD122 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[488] WL[489] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_245 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD122 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[490] WL[491] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS245 DEC_X1_REP[5] SH_NPD122 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_246 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD123 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[492] WL[493] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_247 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[5]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD123 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[494] WL[495] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS247 DEC_X1_REP[5] SH_NPD123 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_248 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD124 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[496] WL[497] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_249 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD124 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[498] WL[499] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS249 DEC_X1_REP[6] SH_NPD124 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_250 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD125 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[500] WL[501] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_251 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[6]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD125 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[502] WL[503] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS251 DEC_X1_REP[6] SH_NPD125 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_252 DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD126 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[504] WL[505] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_253 DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD126 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[506] WL[507] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS253 DEC_X1_REP[7] SH_NPD126 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_254 DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD127 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[508] WL[509] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_255 DEC_X0_REP[6] DEC_X0_REP[7] DEC_X0_REP[0] DEC_X0_REP[1]
+ DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5] DEC_X1_REP[7]
+ DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4]
+ DEC_X1_REP[5] DEC_X1_REP[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SH_NPD127 SLP_LCTRL_REP TK VXDDHD VDDI VSSI WE WL[510] WL[511] WLPY_UP[3]
+ WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS255 DEC_X1_REP[7] SH_NPD127 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_BANK_F_REP GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6]
+ GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15]
+ GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23]
+ GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31]
+ GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6]
+ GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17]
+ GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28]
+ GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3]
+ GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13]
+ GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22]
+ GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31]
+ GWB[32] GWB[33] GWB[34] GWB[35] DSLP_BUF SLP_LCTRL RE WE VXDDHD WLP_SAE
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5]
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1]
+ DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] YL[1] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] VXDDAI
+ VDDI VSSI WLP_SAE_TK TK
XLIO_MCB_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] VXDDAI LIOPD WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7]
+ WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18]
+ WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29]
+ WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40]
+ WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51]
+ WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62]
+ WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73]
+ WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84]
+ WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95]
+ WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105]
+ WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114]
+ WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123]
+ WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] WL[132]
+ WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141]
+ WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150]
+ WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159]
+ WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168]
+ WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177]
+ WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186]
+ WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] WL[195]
+ WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204]
+ WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213]
+ WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222]
+ WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231]
+ WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240]
+ WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249]
+ WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] WL[258]
+ WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] WL[267]
+ WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] WL[276]
+ WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] WL[285]
+ WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] WL[294]
+ WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] WL[303]
+ WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] WL[312]
+ WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] WL[321]
+ WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] WL[330]
+ WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] WL[339]
+ WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] WL[348]
+ WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] WL[357]
+ WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] WL[366]
+ WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] WL[375]
+ WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] WL[383] WL[384]
+ WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] WL[392] WL[393]
+ WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] WL[401] WL[402]
+ WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] WL[410] WL[411]
+ WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] WL[419] WL[420]
+ WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] WL[428] WL[429]
+ WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] WL[437] WL[438]
+ WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] WL[446] WL[447]
+ WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] WL[455] WL[456]
+ WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] WL[464] WL[465]
+ WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] WL[473] WL[474]
+ WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] WL[482] WL[483]
+ WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] WL[491] WL[492]
+ WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] WL[500] WL[501]
+ WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] WL[509] WL[510]
+ WL[511] BLEQ_DN BLEQ_UP GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8]
+ GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19]
+ GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30]
+ GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5]
+ GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15]
+ GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24]
+ GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33]
+ GWB[34] GWB[35] RE_LIO SAEB WE_LIO DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2]
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0]
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6]
+ DEC_Y_UP[7] YL_LIO[0] YL_LIO[1] VDDI VSSI S1BSVTSWSO8000Y24_LIO_MCB_F
XLCTRL_S_M16_SD BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1]
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4]
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4]
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3]
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1]
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7]
+ DSLP_BUF LIOPD RE RE_LIO SAEB SLP_LCTRL TK VXDDHD VDDI VSSI WE WE_LIO
+ WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2]
+ WLPY_UP[3] WLP_SAE WLP_SAE_TK YL[0] YL[1] YL_LIO[0] YL_LIO[1]
+ S1BSVTSWSO8000Y24_LCTRL_S_M16_SD
XXDRV_STRAPD0 VXDDHD VDDI VSSI WLPY_DN[0] WLPY_DNB[0]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_NOR_SHA_0 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD0 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[0]
+ WL[1] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_1 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD0 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[2]
+ WL[3] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS1 DEC_X1[0] SH_NPD0 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_2 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD1 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[4]
+ WL[5] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_3 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD1 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[6]
+ WL[7] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS3 DEC_X1[0] SH_NPD1 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_4 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD2 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[8]
+ WL[9] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_5 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD2 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[10]
+ WL[11] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS5 DEC_X1[1] SH_NPD2 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_6 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD3 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[12]
+ WL[13] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_7 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD3 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[14]
+ WL[15] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS7 DEC_X1[1] SH_NPD3 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_8 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD4 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[16]
+ WL[17] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_9 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD4 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[18]
+ WL[19] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS9 DEC_X1[2] SH_NPD4 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_10 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD5 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[20]
+ WL[21] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_11 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD5 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[22]
+ WL[23] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS11 DEC_X1[2] SH_NPD5 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_12 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD6 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[24]
+ WL[25] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_13 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD6 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[26]
+ WL[27] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS13 DEC_X1[3] SH_NPD6 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_14 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD7 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[28]
+ WL[29] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_15 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD7 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[30]
+ WL[31] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS15 DEC_X1[3] SH_NPD7 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_16 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD8 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[32]
+ WL[33] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_17 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD8 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[34]
+ WL[35] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS17 DEC_X1[4] SH_NPD8 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_18 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD9 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[36]
+ WL[37] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_19 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD9 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[38]
+ WL[39] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS19 DEC_X1[4] SH_NPD9 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_20 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD10 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[40]
+ WL[41] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_21 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD10 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[42]
+ WL[43] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS21 DEC_X1[5] SH_NPD10 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_22 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD11 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[44]
+ WL[45] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_23 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD11 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[46]
+ WL[47] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS23 DEC_X1[5] SH_NPD11 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_24 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD12 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[48]
+ WL[49] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_25 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD12 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[50]
+ WL[51] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS25 DEC_X1[6] SH_NPD12 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_26 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD13 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[52]
+ WL[53] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_27 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD13 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[54]
+ WL[55] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS27 DEC_X1[6] SH_NPD13 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_28 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD14 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[56]
+ WL[57] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_29 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD14 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[58]
+ WL[59] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS29 DEC_X1[7] SH_NPD14 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_30 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD15 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[60]
+ WL[61] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_31 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD15 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[62]
+ WL[63] WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS31 DEC_X1[7] SH_NPD15 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_STRAPD1 VXDDHD VDDI VSSI WLPY_DN[1] WLPY_DNB[1]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_NOR_SHA_32 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD16 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[64]
+ WL[65] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_33 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD16 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[66]
+ WL[67] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS33 DEC_X1[0] SH_NPD16 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_34 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD17 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[68]
+ WL[69] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_35 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD17 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[70]
+ WL[71] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS35 DEC_X1[0] SH_NPD17 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_36 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD18 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[72]
+ WL[73] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_37 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD18 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[74]
+ WL[75] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS37 DEC_X1[1] SH_NPD18 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_38 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD19 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[76]
+ WL[77] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_39 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD19 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[78]
+ WL[79] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS39 DEC_X1[1] SH_NPD19 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_40 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD20 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[80]
+ WL[81] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_41 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD20 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[82]
+ WL[83] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS41 DEC_X1[2] SH_NPD20 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_42 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD21 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[84]
+ WL[85] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_43 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD21 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[86]
+ WL[87] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS43 DEC_X1[2] SH_NPD21 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_44 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD22 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[88]
+ WL[89] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_45 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD22 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[90]
+ WL[91] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS45 DEC_X1[3] SH_NPD22 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_46 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD23 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[92]
+ WL[93] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_47 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD23 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[94]
+ WL[95] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS47 DEC_X1[3] SH_NPD23 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_48 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD24 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[96]
+ WL[97] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_49 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD24 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[98]
+ WL[99] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS49 DEC_X1[4] SH_NPD24 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_50 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD25 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[100] WL[101] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_51 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD25 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[102] WL[103] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS51 DEC_X1[4] SH_NPD25 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_52 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD26 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[104] WL[105] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_53 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD26 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[106] WL[107] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS53 DEC_X1[5] SH_NPD26 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_54 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD27 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[108] WL[109] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_55 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD27 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[110] WL[111] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS55 DEC_X1[5] SH_NPD27 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_56 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD28 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[112] WL[113] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_57 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD28 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[114] WL[115] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS57 DEC_X1[6] SH_NPD28 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_58 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD29 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[116] WL[117] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_59 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD29 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[118] WL[119] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS59 DEC_X1[6] SH_NPD29 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_60 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD30 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[120] WL[121] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_61 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD30 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[122] WL[123] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS61 DEC_X1[7] SH_NPD30 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_62 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD31 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[124] WL[125] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_63 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD31 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[126] WL[127] WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS63 DEC_X1[7] SH_NPD31 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_STRAPD2 VXDDHD VDDI VSSI WLPY_DN[2] WLPY_DNB[2]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_NOR_SHA_64 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD32 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[128] WL[129] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_65 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD32 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[130] WL[131] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS65 DEC_X1[0] SH_NPD32 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_66 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD33 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[132] WL[133] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_67 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD33 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[134] WL[135] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS67 DEC_X1[0] SH_NPD33 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_68 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD34 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[136] WL[137] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_69 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD34 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[138] WL[139] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS69 DEC_X1[1] SH_NPD34 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_70 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD35 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[140] WL[141] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_71 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD35 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[142] WL[143] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS71 DEC_X1[1] SH_NPD35 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_72 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD36 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[144] WL[145] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_73 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD36 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[146] WL[147] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS73 DEC_X1[2] SH_NPD36 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_74 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD37 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[148] WL[149] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_75 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD37 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[150] WL[151] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS75 DEC_X1[2] SH_NPD37 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_76 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD38 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[152] WL[153] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_77 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD38 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[154] WL[155] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS77 DEC_X1[3] SH_NPD38 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_78 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD39 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[156] WL[157] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_79 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD39 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[158] WL[159] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS79 DEC_X1[3] SH_NPD39 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_80 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD40 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[160] WL[161] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_81 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD40 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[162] WL[163] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS81 DEC_X1[4] SH_NPD40 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_82 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD41 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[164] WL[165] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_83 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD41 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[166] WL[167] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS83 DEC_X1[4] SH_NPD41 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_84 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD42 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[168] WL[169] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_85 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD42 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[170] WL[171] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS85 DEC_X1[5] SH_NPD42 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_86 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD43 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[172] WL[173] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_87 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD43 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[174] WL[175] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS87 DEC_X1[5] SH_NPD43 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_88 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD44 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[176] WL[177] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_89 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD44 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[178] WL[179] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS89 DEC_X1[6] SH_NPD44 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_90 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD45 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[180] WL[181] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_91 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD45 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[182] WL[183] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS91 DEC_X1[6] SH_NPD45 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_92 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD46 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[184] WL[185] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_93 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD46 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[186] WL[187] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS93 DEC_X1[7] SH_NPD46 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_94 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD47 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[188] WL[189] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_95 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD47 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[190] WL[191] WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS95 DEC_X1[7] SH_NPD47 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_STRAPD3 VXDDHD VDDI VSSI WLPY_DN[3] WLPY_DNB[3]
+ S1BSVTSWSO8000Y24_XDRV_STRAP_LCNT
XXDRV_LA512_NOR_SHA_96 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD48 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[192] WL[193] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_97 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD48 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[194] WL[195] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS97 DEC_X1[0] SH_NPD48 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_98 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD49 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[196] WL[197] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_99 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD49 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[198] WL[199] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS99 DEC_X1[0] SH_NPD49 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_100 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD50 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[200] WL[201] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_101 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD50 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[202] WL[203] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS101 DEC_X1[1] SH_NPD50 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_102 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD51 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[204] WL[205] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_103 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD51 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[206] WL[207] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS103 DEC_X1[1] SH_NPD51 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_104 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD52 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[208] WL[209] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_105 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD52 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[210] WL[211] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS105 DEC_X1[2] SH_NPD52 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_106 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD53 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[212] WL[213] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_107 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD53 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[214] WL[215] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS107 DEC_X1[2] SH_NPD53 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_108 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD54 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[216] WL[217] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_109 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD54 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[218] WL[219] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS109 DEC_X1[3] SH_NPD54 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_110 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD55 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[220] WL[221] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_111 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD55 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[222] WL[223] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS111 DEC_X1[3] SH_NPD55 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_112 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD56 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[224] WL[225] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_113 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD56 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[226] WL[227] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS113 DEC_X1[4] SH_NPD56 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_114 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD57 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[228] WL[229] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_115 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD57 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[230] WL[231] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS115 DEC_X1[4] SH_NPD57 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_116 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD58 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[232] WL[233] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_117 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD58 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[234] WL[235] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS117 DEC_X1[5] SH_NPD58 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_118 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD59 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[236] WL[237] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_119 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD59 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[238] WL[239] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS119 DEC_X1[5] SH_NPD59 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_120 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD60 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[240] WL[241] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_121 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD60 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[242] WL[243] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS121 DEC_X1[6] SH_NPD60 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_122 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD61 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[244] WL[245] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_123 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD61 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[246] WL[247] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS123 DEC_X1[6] SH_NPD61 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_124 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD62 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[248] WL[249] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_125 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD62 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[250] WL[251] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS125 DEC_X1[7] SH_NPD62 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_126 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD63 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[252] WL[253] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_127 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD63 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[254] WL[255] WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS127 DEC_X1[7] SH_NPD63 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_STRAPU0 VXDDHD VDDI VSSI WLPY_UP[0] WLPY_UPB[0]
+ S1BSVTSWSO8000Y24_XDRV_STRAP_LCNT
XXDRV_LA512_NOR_SHA_128 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD64 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[256] WL[257] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_129 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD64 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[258] WL[259] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS129 DEC_X1[0] SH_NPD64 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_130 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD65 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[260] WL[261] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_131 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD65 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[262] WL[263] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS131 DEC_X1[0] SH_NPD65 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_132 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD66 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[264] WL[265] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_133 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD66 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[266] WL[267] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS133 DEC_X1[1] SH_NPD66 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_134 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD67 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[268] WL[269] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_135 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD67 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[270] WL[271] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS135 DEC_X1[1] SH_NPD67 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_136 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD68 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[272] WL[273] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_137 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD68 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[274] WL[275] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS137 DEC_X1[2] SH_NPD68 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_138 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD69 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[276] WL[277] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_139 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD69 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[278] WL[279] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS139 DEC_X1[2] SH_NPD69 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_140 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD70 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[280] WL[281] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_141 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD70 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[282] WL[283] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS141 DEC_X1[3] SH_NPD70 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_142 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD71 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[284] WL[285] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_143 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD71 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[286] WL[287] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS143 DEC_X1[3] SH_NPD71 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_144 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD72 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[288] WL[289] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_145 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD72 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[290] WL[291] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS145 DEC_X1[4] SH_NPD72 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_146 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD73 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[292] WL[293] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_147 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD73 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[294] WL[295] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS147 DEC_X1[4] SH_NPD73 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_148 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD74 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[296] WL[297] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_149 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD74 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[298] WL[299] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS149 DEC_X1[5] SH_NPD74 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_150 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD75 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[300] WL[301] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_151 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD75 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[302] WL[303] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS151 DEC_X1[5] SH_NPD75 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_152 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD76 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[304] WL[305] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_153 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD76 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[306] WL[307] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS153 DEC_X1[6] SH_NPD76 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_154 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD77 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[308] WL[309] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_155 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD77 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[310] WL[311] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS155 DEC_X1[6] SH_NPD77 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_156 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD78 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[312] WL[313] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_157 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD78 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[314] WL[315] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS157 DEC_X1[7] SH_NPD78 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_158 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD79 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[316] WL[317] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_159 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD79 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[318] WL[319] WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS159 DEC_X1[7] SH_NPD79 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_STRAPU1 VXDDHD VDDI VSSI WLPY_UP[1] WLPY_UPB[1]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_NOR_SHA_160 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD80 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[320] WL[321] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_161 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD80 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[322] WL[323] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS161 DEC_X1[0] SH_NPD80 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_162 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD81 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[324] WL[325] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_163 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD81 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[326] WL[327] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS163 DEC_X1[0] SH_NPD81 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_164 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD82 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[328] WL[329] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_165 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD82 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[330] WL[331] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS165 DEC_X1[1] SH_NPD82 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_166 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD83 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[332] WL[333] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_167 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD83 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[334] WL[335] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS167 DEC_X1[1] SH_NPD83 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_168 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD84 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[336] WL[337] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_169 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD84 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[338] WL[339] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS169 DEC_X1[2] SH_NPD84 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_170 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD85 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[340] WL[341] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_171 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD85 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[342] WL[343] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS171 DEC_X1[2] SH_NPD85 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_172 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD86 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[344] WL[345] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_173 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD86 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[346] WL[347] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS173 DEC_X1[3] SH_NPD86 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_174 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD87 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[348] WL[349] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_175 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD87 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[350] WL[351] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS175 DEC_X1[3] SH_NPD87 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_176 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD88 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[352] WL[353] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_177 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD88 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[354] WL[355] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS177 DEC_X1[4] SH_NPD88 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_178 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD89 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[356] WL[357] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_179 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD89 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[358] WL[359] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS179 DEC_X1[4] SH_NPD89 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_180 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD90 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[360] WL[361] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_181 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD90 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[362] WL[363] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS181 DEC_X1[5] SH_NPD90 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_182 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD91 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[364] WL[365] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_183 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD91 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[366] WL[367] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS183 DEC_X1[5] SH_NPD91 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_184 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD92 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[368] WL[369] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_185 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD92 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[370] WL[371] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS185 DEC_X1[6] SH_NPD92 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_186 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD93 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[372] WL[373] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_187 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD93 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[374] WL[375] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS187 DEC_X1[6] SH_NPD93 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_188 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD94 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[376] WL[377] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_189 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD94 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[378] WL[379] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS189 DEC_X1[7] SH_NPD94 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_190 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD95 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[380] WL[381] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_191 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD95 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[382] WL[383] WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS191 DEC_X1[7] SH_NPD95 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_STRAPU2 VXDDHD VDDI VSSI WLPY_UP[2] WLPY_UPB[2]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_NOR_SHA_192 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD96 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[384] WL[385] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_193 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD96 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[386] WL[387] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS193 DEC_X1[0] SH_NPD96 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_194 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD97 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[388] WL[389] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_195 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD97 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[390] WL[391] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS195 DEC_X1[0] SH_NPD97 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_196 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD98 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[392] WL[393] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_197 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD98 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[394] WL[395] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS197 DEC_X1[1] SH_NPD98 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_198 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD99 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[396] WL[397] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_199 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD99 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[398] WL[399] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS199 DEC_X1[1] SH_NPD99 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_200 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD100 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[400] WL[401] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_201 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD100 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[402] WL[403] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS201 DEC_X1[2] SH_NPD100 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_202 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD101 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[404] WL[405] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_203 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD101 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[406] WL[407] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS203 DEC_X1[2] SH_NPD101 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_204 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD102 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[408] WL[409] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_205 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD102 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[410] WL[411] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS205 DEC_X1[3] SH_NPD102 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_206 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD103 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[412] WL[413] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_207 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD103 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[414] WL[415] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS207 DEC_X1[3] SH_NPD103 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_208 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD104 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[416] WL[417] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_209 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD104 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[418] WL[419] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS209 DEC_X1[4] SH_NPD104 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_210 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD105 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[420] WL[421] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_211 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD105 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[422] WL[423] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS211 DEC_X1[4] SH_NPD105 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_212 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD106 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[424] WL[425] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_213 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD106 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[426] WL[427] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS213 DEC_X1[5] SH_NPD106 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_214 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD107 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[428] WL[429] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_215 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD107 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[430] WL[431] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS215 DEC_X1[5] SH_NPD107 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_216 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD108 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[432] WL[433] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_217 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD108 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[434] WL[435] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS217 DEC_X1[6] SH_NPD108 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_218 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD109 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[436] WL[437] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_219 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD109 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[438] WL[439] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS219 DEC_X1[6] SH_NPD109 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_220 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD110 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[440] WL[441] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_221 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD110 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[442] WL[443] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS221 DEC_X1[7] SH_NPD110 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_222 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD111 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[444] WL[445] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_223 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD111 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[446] WL[447] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS223 DEC_X1[7] SH_NPD111 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_STRAPU3 VXDDHD VDDI VSSI WLPY_UP[3] WLPY_UPB[3]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_NOR_SHA_224 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD112 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[448] WL[449] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_225 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD112 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[450] WL[451] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS225 DEC_X1[0] SH_NPD112 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_226 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD113 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[452] WL[453] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_227 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD113 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[454] WL[455] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS227 DEC_X1[0] SH_NPD113 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_228 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD114 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[456] WL[457] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_229 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD114 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[458] WL[459] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS229 DEC_X1[1] SH_NPD114 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_230 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD115 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[460] WL[461] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_231 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD115 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[462] WL[463] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS231 DEC_X1[1] SH_NPD115 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_232 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD116 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[464] WL[465] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_233 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD116 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[466] WL[467] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS233 DEC_X1[2] SH_NPD116 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_234 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD117 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[468] WL[469] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_235 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD117 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[470] WL[471] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS235 DEC_X1[2] SH_NPD117 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_236 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD118 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[472] WL[473] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_237 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD118 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[474] WL[475] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS237 DEC_X1[3] SH_NPD118 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_238 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD119 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[476] WL[477] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_239 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD119 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[478] WL[479] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS239 DEC_X1[3] SH_NPD119 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_240 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD120 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[480] WL[481] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_241 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD120 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[482] WL[483] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS241 DEC_X1[4] SH_NPD120 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_242 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD121 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[484] WL[485] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_243 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD121 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[486] WL[487] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS243 DEC_X1[4] SH_NPD121 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_244 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD122 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[488] WL[489] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_245 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD122 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[490] WL[491] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS245 DEC_X1[5] SH_NPD122 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_246 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD123 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[492] WL[493] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_247 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD123 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[494] WL[495] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS247 DEC_X1[5] SH_NPD123 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_248 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD124 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[496] WL[497] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_249 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD124 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[498] WL[499] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS249 DEC_X1[6] SH_NPD124 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_250 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD125 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[500] WL[501] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_251 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD125 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[502] WL[503] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS251 DEC_X1[6] SH_NPD125 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_252 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD126 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[504] WL[505] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_253 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD126 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[506] WL[507] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS253 DEC_X1[7] SH_NPD126 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
XXDRV_LA512_NOR_SHA_254 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD127 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[508] WL[509] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_NOR_SHA_255 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DSLP_BUF RE SH_NPD127 SLP_LCTRL TK VXDDHD VDDI VSSI WE
+ WL[510] WL[511] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_NOR_SHA
XXDRV_LA512_SHA_PMOS255 DEC_X1[7] SH_NPD127 VDDI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_PMOS
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_WL_TRK WL_TK BL_TK SLP_BUF VXDDHD TIEH TIEL VXDDAI
+ VDDI VSSI
XTKWL_2X2_RL0 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL1 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL2 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL3 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL4 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL5 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL6 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL7 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL8 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL9 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL10 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL11 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL12 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL13 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL14 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL15 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL16 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL17 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL18 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL19 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL20 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL21 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL22 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL23 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL24 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL25 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL26 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL27 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL28 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL29 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL30 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL31 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL32 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL33 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL34 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL35 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL36 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL37 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL38 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL39 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL40 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL41 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL42 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL43 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL44 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL45 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL46 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL47 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL48 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL49 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL50 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL51 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL52 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL53 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL54 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL55 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL56 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL57 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL58 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL59 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL60 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL61 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL62 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL63 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL64 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL65 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL66 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL67 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL68 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL69 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL70 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL71 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RL72 VXDDAI VDDI VSSI WL_TK WL_TK S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_ISO VXDDAI VDDI VSSI WL_TK WL_TK TIEL TIEL
+ S1BSVTSWSO8000Y24_TKWL_2X2_ISO
XTKWL_2X2_RR0 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR1 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR2 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR3 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR4 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR5 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR6 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR7 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR8 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR9 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR10 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR11 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR12 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR13 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR14 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR15 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR16 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR17 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR18 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR19 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR20 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR21 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR22 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR23 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR24 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR25 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR26 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR27 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR28 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR29 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR30 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR31 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR32 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR33 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR34 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR35 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR36 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR37 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR38 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR39 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR40 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR41 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR42 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR43 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR44 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR45 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR46 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR47 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR48 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR49 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR50 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR51 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR52 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR53 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR54 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR55 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR56 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR57 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR58 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR59 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR60 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR61 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR62 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR63 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR64 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR65 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR66 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR67 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR68 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR69 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_RR70 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKBL_TRKPRE SLP_BUF BL_TK WL_TK VXDDAI VDDI VSSI TIEH TIEL
+ S1BSVTSWSO8000Y24_TKBL_TRKPRE
XTKWL_2X2_L0 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L1 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L2 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L3 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L4 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L5 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L6 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L7 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L8 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L9 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L10 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L11 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L12 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L13 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L14 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L15 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L16 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L17 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L18 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L19 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L20 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L21 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L22 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L23 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L24 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L25 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L26 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L27 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L28 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L29 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L30 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L31 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L32 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L33 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L34 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L35 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L36 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L37 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L38 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L39 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L40 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L41 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L42 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L43 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L44 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L45 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L46 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L47 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L48 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L49 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L50 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L51 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L52 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L53 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L54 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L55 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L56 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L57 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L58 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L59 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L60 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L61 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L62 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L63 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L64 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L65 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L66 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L67 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L68 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L69 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L70 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L71 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L72 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L73 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L74 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L75 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L76 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L77 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L78 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L79 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L80 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L81 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L82 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L83 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L84 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L85 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L86 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L87 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L88 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L89 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L90 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L91 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L92 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L93 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L94 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L95 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L96 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L97 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L98 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L99 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L100 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L101 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L102 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L103 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L104 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L105 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L106 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L107 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L108 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L109 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L110 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L111 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L112 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L113 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L114 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L115 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L116 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L117 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L118 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L119 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L120 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L121 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L122 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L123 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L124 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L125 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L126 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L127 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L128 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L129 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L130 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L131 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L132 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L133 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L134 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L135 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L136 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L137 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L138 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L139 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L140 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L141 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L142 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
XTKWL_2X2_L143 VXDDAI VDDI VSSI TIEL TIEL S1BSVTSWSO8000Y24_TKWL_2X2
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_TRACKING WL_TK SLP_BUF BL_TK VXDDHD WL[0] WL[1] WL[2]
+ WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14]
+ WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25]
+ WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36]
+ WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47]
+ WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58]
+ WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69]
+ WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80]
+ WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91]
+ WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101]
+ WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110]
+ WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119]
+ WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128]
+ WL[129] WL[130] WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137]
+ WL[138] WL[139] WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146]
+ WL[147] WL[148] WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155]
+ WL[156] WL[157] WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164]
+ WL[165] WL[166] WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173]
+ WL[174] WL[175] WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182]
+ WL[183] WL[184] WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191]
+ WL[192] WL[193] WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200]
+ WL[201] WL[202] WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209]
+ WL[210] WL[211] WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218]
+ WL[219] WL[220] WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227]
+ WL[228] WL[229] WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236]
+ WL[237] WL[238] WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245]
+ WL[246] WL[247] WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254]
+ WL[255] VXDDAI VDDI VSSI
XWL_TRK WL_TK BL_TK SLP_BUF VXDDHD TIEH TIEL VXDDAI VDDI VSSI
+ S1BSVTSWSO8000Y24_WL_TRK
X0TRKNORX2_0 BL_TK VXDDAI VDDI VSSI WL[0] WL[1] WL_TK FLOAT1[0] NET[0] FLOAT3
+ NET_TRKBL[0] FLOAT5 TIEH S1BSVTSWSO8000Y24_TRKNORX2
X1TRKNORX2_1 BL_TK VXDDAI VDDI VSSI WL[2] WL[3] WL_TK FLOAT1[1] NET[1] NET[0]
+ NET_TRKBL[1] NET_TRKBL[0] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X2TRKNORX2_2 BL_TK VXDDAI VDDI VSSI WL[4] WL[5] WL_TK FLOAT1[2] NET[2] NET[1]
+ NET_TRKBL[2] NET_TRKBL[1] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X3TRKNORX2_3 BL_TK VXDDAI VDDI VSSI WL[6] WL[7] WL_TK FLOAT1[3] NET[3] NET[2]
+ NET_TRKBL[3] NET_TRKBL[2] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_4 BL_TK VXDDAI VDDI VSSI WL[8] WL[9] TIEL FLOAT1[4] NET[4] NET[3]
+ NET_TRKBL[4] NET_TRKBL[3] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_5 BL_TK VXDDAI VDDI VSSI WL[10] WL[11] TIEL FLOAT1[5] NET[5] NET[4]
+ NET_TRKBL[5] NET_TRKBL[4] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_6 BL_TK VXDDAI VDDI VSSI WL[12] WL[13] TIEL FLOAT1[6] NET[6] NET[5]
+ NET_TRKBL[6] NET_TRKBL[5] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_7 BL_TK VXDDAI VDDI VSSI WL[14] WL[15] TIEL FLOAT1[7] NET[7] NET[6]
+ NET_TRKBL[7] NET_TRKBL[6] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_8 BL_TK VXDDAI VDDI VSSI WL[16] WL[17] TIEL FLOAT1[8] NET[8] NET[7]
+ NET_TRKBL[8] NET_TRKBL[7] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_9 BL_TK VXDDAI VDDI VSSI WL[18] WL[19] TIEL FLOAT1[9] NET[9] NET[8]
+ NET_TRKBL[9] NET_TRKBL[8] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_10 BL_TK VXDDAI VDDI VSSI WL[20] WL[21] TIEL FLOAT1[10] NET[10]
+ NET[9] NET_TRKBL[10] NET_TRKBL[9] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_11 BL_TK VXDDAI VDDI VSSI WL[22] WL[23] TIEL FLOAT1[11] NET[11]
+ NET[10] NET_TRKBL[11] NET_TRKBL[10] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_12 BL_TK VXDDAI VDDI VSSI WL[24] WL[25] TIEL FLOAT1[12] NET[12]
+ NET[11] NET_TRKBL[12] NET_TRKBL[11] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_13 BL_TK VXDDAI VDDI VSSI WL[26] WL[27] TIEL FLOAT1[13] NET[13]
+ NET[12] NET_TRKBL[13] NET_TRKBL[12] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_14 BL_TK VXDDAI VDDI VSSI WL[28] WL[29] TIEL FLOAT1[14] NET[14]
+ NET[13] NET_TRKBL[14] NET_TRKBL[13] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_15 BL_TK VXDDAI VDDI VSSI WL[30] WL[31] TIEL FLOAT1[15] NET[15]
+ NET[14] NET_TRKBL[15] NET_TRKBL[14] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_16 BL_TK VXDDAI VDDI VSSI WL[32] WL[33] TIEL FLOAT1[16] NET[16]
+ NET[15] NET_TRKBL[16] NET_TRKBL[15] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_17 BL_TK VXDDAI VDDI VSSI WL[34] WL[35] TIEL FLOAT1[17] NET[17]
+ NET[16] NET_TRKBL[17] NET_TRKBL[16] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_18 BL_TK VXDDAI VDDI VSSI WL[36] WL[37] TIEL FLOAT1[18] NET[18]
+ NET[17] NET_TRKBL[18] NET_TRKBL[17] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_19 BL_TK VXDDAI VDDI VSSI WL[38] WL[39] TIEL FLOAT1[19] NET[19]
+ NET[18] NET_TRKBL[19] NET_TRKBL[18] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_20 BL_TK VXDDAI VDDI VSSI WL[40] WL[41] TIEL FLOAT1[20] NET[20]
+ NET[19] NET_TRKBL[20] NET_TRKBL[19] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_21 BL_TK VXDDAI VDDI VSSI WL[42] WL[43] TIEL FLOAT1[21] NET[21]
+ NET[20] NET_TRKBL[21] NET_TRKBL[20] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_22 BL_TK VXDDAI VDDI VSSI WL[44] WL[45] TIEL FLOAT1[22] NET[22]
+ NET[21] NET_TRKBL[22] NET_TRKBL[21] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_23 BL_TK VXDDAI VDDI VSSI WL[46] WL[47] TIEL FLOAT1[23] NET[23]
+ NET[22] NET_TRKBL[23] NET_TRKBL[22] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_24 BL_TK VXDDAI VDDI VSSI WL[48] WL[49] TIEL FLOAT1[24] NET[24]
+ NET[23] NET_TRKBL[24] NET_TRKBL[23] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_25 BL_TK VXDDAI VDDI VSSI WL[50] WL[51] TIEL FLOAT1[25] NET[25]
+ NET[24] NET_TRKBL[25] NET_TRKBL[24] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_26 BL_TK VXDDAI VDDI VSSI WL[52] WL[53] TIEL FLOAT1[26] NET[26]
+ NET[25] NET_TRKBL[26] NET_TRKBL[25] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_27 BL_TK VXDDAI VDDI VSSI WL[54] WL[55] TIEL FLOAT1[27] NET[27]
+ NET[26] NET_TRKBL[27] NET_TRKBL[26] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_28 BL_TK VXDDAI VDDI VSSI WL[56] WL[57] TIEL FLOAT1[28] NET[28]
+ NET[27] NET_TRKBL[28] NET_TRKBL[27] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_29 BL_TK VXDDAI VDDI VSSI WL[58] WL[59] TIEL FLOAT1[29] NET[29]
+ NET[28] NET_TRKBL[29] NET_TRKBL[28] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_30 BL_TK VXDDAI VDDI VSSI WL[60] WL[61] TIEL FLOAT1[30] NET[30]
+ NET[29] NET_TRKBL[30] NET_TRKBL[29] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_31 BL_TK VXDDAI VDDI VSSI WL[62] WL[63] TIEL FLOAT1[31] NET[31]
+ NET[30] NET_TRKBL[31] NET_TRKBL[30] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_32 BL_TK VXDDAI VDDI VSSI WL[64] WL[65] TIEL FLOAT1[32] NET[32]
+ NET[31] NET_TRKBL[32] NET_TRKBL[31] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_33 BL_TK VXDDAI VDDI VSSI WL[66] WL[67] TIEL FLOAT1[33] NET[33]
+ NET[32] NET_TRKBL[33] NET_TRKBL[32] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_34 BL_TK VXDDAI VDDI VSSI WL[68] WL[69] TIEL FLOAT1[34] NET[34]
+ NET[33] NET_TRKBL[34] NET_TRKBL[33] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_35 BL_TK VXDDAI VDDI VSSI WL[70] WL[71] TIEL FLOAT1[35] NET[35]
+ NET[34] NET_TRKBL[35] NET_TRKBL[34] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_36 BL_TK VXDDAI VDDI VSSI WL[72] WL[73] TIEL FLOAT1[36] NET[36]
+ NET[35] NET_TRKBL[36] NET_TRKBL[35] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_37 BL_TK VXDDAI VDDI VSSI WL[74] WL[75] TIEL FLOAT1[37] NET[37]
+ NET[36] NET_TRKBL[37] NET_TRKBL[36] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_38 BL_TK VXDDAI VDDI VSSI WL[76] WL[77] TIEL FLOAT1[38] NET[38]
+ NET[37] NET_TRKBL[38] NET_TRKBL[37] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_39 BL_TK VXDDAI VDDI VSSI WL[78] WL[79] TIEL FLOAT1[39] NET[39]
+ NET[38] NET_TRKBL[39] NET_TRKBL[38] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_40 BL_TK VXDDAI VDDI VSSI WL[80] WL[81] TIEL FLOAT1[40] NET[40]
+ NET[39] NET_TRKBL[40] NET_TRKBL[39] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_41 BL_TK VXDDAI VDDI VSSI WL[82] WL[83] TIEL FLOAT1[41] NET[41]
+ NET[40] NET_TRKBL[41] NET_TRKBL[40] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_42 BL_TK VXDDAI VDDI VSSI WL[84] WL[85] TIEL FLOAT1[42] NET[42]
+ NET[41] NET_TRKBL[42] NET_TRKBL[41] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_43 BL_TK VXDDAI VDDI VSSI WL[86] WL[87] TIEL FLOAT1[43] NET[43]
+ NET[42] NET_TRKBL[43] NET_TRKBL[42] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_44 BL_TK VXDDAI VDDI VSSI WL[88] WL[89] TIEL FLOAT1[44] NET[44]
+ NET[43] NET_TRKBL[44] NET_TRKBL[43] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_45 BL_TK VXDDAI VDDI VSSI WL[90] WL[91] TIEL FLOAT1[45] NET[45]
+ NET[44] NET_TRKBL[45] NET_TRKBL[44] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_46 BL_TK VXDDAI VDDI VSSI WL[92] WL[93] TIEL FLOAT1[46] NET[46]
+ NET[45] NET_TRKBL[46] NET_TRKBL[45] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_47 BL_TK VXDDAI VDDI VSSI WL[94] WL[95] TIEL FLOAT1[47] NET[47]
+ NET[46] NET_TRKBL[47] NET_TRKBL[46] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_48 BL_TK VXDDAI VDDI VSSI WL[96] WL[97] TIEL FLOAT1[48] NET[48]
+ NET[47] NET_TRKBL[48] NET_TRKBL[47] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_49 BL_TK VXDDAI VDDI VSSI WL[98] WL[99] TIEL FLOAT1[49] NET[49]
+ NET[48] NET_TRKBL[49] NET_TRKBL[48] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_50 BL_TK VXDDAI VDDI VSSI WL[100] WL[101] TIEL FLOAT1[50] NET[50]
+ NET[49] NET_TRKBL[50] NET_TRKBL[49] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_51 BL_TK VXDDAI VDDI VSSI WL[102] WL[103] TIEL FLOAT1[51] NET[51]
+ NET[50] NET_TRKBL[51] NET_TRKBL[50] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_52 BL_TK VXDDAI VDDI VSSI WL[104] WL[105] TIEL FLOAT1[52] NET[52]
+ NET[51] NET_TRKBL[52] NET_TRKBL[51] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_53 BL_TK VXDDAI VDDI VSSI WL[106] WL[107] TIEL FLOAT1[53] NET[53]
+ NET[52] NET_TRKBL[53] NET_TRKBL[52] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_54 BL_TK VXDDAI VDDI VSSI WL[108] WL[109] TIEL FLOAT1[54] NET[54]
+ NET[53] NET_TRKBL[54] NET_TRKBL[53] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_55 BL_TK VXDDAI VDDI VSSI WL[110] WL[111] TIEL FLOAT1[55] NET[55]
+ NET[54] NET_TRKBL[55] NET_TRKBL[54] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_56 BL_TK VXDDAI VDDI VSSI WL[112] WL[113] TIEL FLOAT1[56] NET[56]
+ NET[55] NET_TRKBL[56] NET_TRKBL[55] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_57 BL_TK VXDDAI VDDI VSSI WL[114] WL[115] TIEL FLOAT1[57] NET[57]
+ NET[56] NET_TRKBL[57] NET_TRKBL[56] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_58 BL_TK VXDDAI VDDI VSSI WL[116] WL[117] TIEL FLOAT1[58] NET[58]
+ NET[57] NET_TRKBL[58] NET_TRKBL[57] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_59 BL_TK VXDDAI VDDI VSSI WL[118] WL[119] TIEL FLOAT1[59] NET[59]
+ NET[58] NET_TRKBL[59] NET_TRKBL[58] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_60 BL_TK VXDDAI VDDI VSSI WL[120] WL[121] TIEL FLOAT1[60] NET[60]
+ NET[59] NET_TRKBL[60] NET_TRKBL[59] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_61 BL_TK VXDDAI VDDI VSSI WL[122] WL[123] TIEL FLOAT1[61] NET[61]
+ NET[60] NET_TRKBL[61] NET_TRKBL[60] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_62 BL_TK VXDDAI VDDI VSSI WL[124] WL[125] TIEL FLOAT1[62] NET[62]
+ NET[61] NET_TRKBL[62] NET_TRKBL[61] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_63 BL_TK VXDDAI VDDI VSSI WL[126] WL[127] TIEL FLOAT1[63] NET[63]
+ NET[62] NET_TRKBL[63] NET_TRKBL[62] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X6TRKNORX2_64 BL_TK VXDDAI VDDI VSSI WL[128] WL[129] TIEL FLOAT1[64] NET[64]
+ NETX[63] NET_TRKBL[64] NET_TRKBLX[63] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_65 BL_TK VXDDAI VDDI VSSI WL[130] WL[131] TIEL FLOAT1[65] NET[65]
+ NET[64] NET_TRKBL[65] NET_TRKBL[64] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_66 BL_TK VXDDAI VDDI VSSI WL[132] WL[133] TIEL FLOAT1[66] NET[66]
+ NET[65] NET_TRKBL[66] NET_TRKBL[65] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_67 BL_TK VXDDAI VDDI VSSI WL[134] WL[135] TIEL FLOAT1[67] NET[67]
+ NET[66] NET_TRKBL[67] NET_TRKBL[66] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_68 BL_TK VXDDAI VDDI VSSI WL[136] WL[137] TIEL FLOAT1[68] NET[68]
+ NET[67] NET_TRKBL[68] NET_TRKBL[67] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_69 BL_TK VXDDAI VDDI VSSI WL[138] WL[139] TIEL FLOAT1[69] NET[69]
+ NET[68] NET_TRKBL[69] NET_TRKBL[68] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_70 BL_TK VXDDAI VDDI VSSI WL[140] WL[141] TIEL FLOAT1[70] NET[70]
+ NET[69] NET_TRKBL[70] NET_TRKBL[69] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_71 BL_TK VXDDAI VDDI VSSI WL[142] WL[143] TIEL FLOAT1[71] NET[71]
+ NET[70] NET_TRKBL[71] NET_TRKBL[70] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_72 BL_TK VXDDAI VDDI VSSI WL[144] WL[145] TIEL FLOAT1[72] NET[72]
+ NET[71] NET_TRKBL[72] NET_TRKBL[71] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_73 BL_TK VXDDAI VDDI VSSI WL[146] WL[147] TIEL FLOAT1[73] NET[73]
+ NET[72] NET_TRKBL[73] NET_TRKBL[72] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_74 BL_TK VXDDAI VDDI VSSI WL[148] WL[149] TIEL FLOAT1[74] NET[74]
+ NET[73] NET_TRKBL[74] NET_TRKBL[73] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_75 BL_TK VXDDAI VDDI VSSI WL[150] WL[151] TIEL FLOAT1[75] NET[75]
+ NET[74] NET_TRKBL[75] NET_TRKBL[74] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_76 BL_TK VXDDAI VDDI VSSI WL[152] WL[153] TIEL FLOAT1[76] NET[76]
+ NET[75] NET_TRKBL[76] NET_TRKBL[75] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_77 BL_TK VXDDAI VDDI VSSI WL[154] WL[155] TIEL FLOAT1[77] NET[77]
+ NET[76] NET_TRKBL[77] NET_TRKBL[76] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_78 BL_TK VXDDAI VDDI VSSI WL[156] WL[157] TIEL FLOAT1[78] NET[78]
+ NET[77] NET_TRKBL[78] NET_TRKBL[77] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_79 BL_TK VXDDAI VDDI VSSI WL[158] WL[159] TIEL FLOAT1[79] NET[79]
+ NET[78] NET_TRKBL[79] NET_TRKBL[78] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_80 BL_TK VXDDAI VDDI VSSI WL[160] WL[161] TIEL FLOAT1[80] NET[80]
+ NET[79] NET_TRKBL[80] NET_TRKBL[79] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_81 BL_TK VXDDAI VDDI VSSI WL[162] WL[163] TIEL FLOAT1[81] NET[81]
+ NET[80] NET_TRKBL[81] NET_TRKBL[80] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_82 BL_TK VXDDAI VDDI VSSI WL[164] WL[165] TIEL FLOAT1[82] NET[82]
+ NET[81] NET_TRKBL[82] NET_TRKBL[81] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_83 BL_TK VXDDAI VDDI VSSI WL[166] WL[167] TIEL FLOAT1[83] NET[83]
+ NET[82] NET_TRKBL[83] NET_TRKBL[82] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_84 BL_TK VXDDAI VDDI VSSI WL[168] WL[169] TIEL FLOAT1[84] NET[84]
+ NET[83] NET_TRKBL[84] NET_TRKBL[83] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_85 BL_TK VXDDAI VDDI VSSI WL[170] WL[171] TIEL FLOAT1[85] NET[85]
+ NET[84] NET_TRKBL[85] NET_TRKBL[84] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_86 BL_TK VXDDAI VDDI VSSI WL[172] WL[173] TIEL FLOAT1[86] NET[86]
+ NET[85] NET_TRKBL[86] NET_TRKBL[85] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_87 BL_TK VXDDAI VDDI VSSI WL[174] WL[175] TIEL FLOAT1[87] NET[87]
+ NET[86] NET_TRKBL[87] NET_TRKBL[86] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_88 BL_TK VXDDAI VDDI VSSI WL[176] WL[177] TIEL FLOAT1[88] NET[88]
+ NET[87] NET_TRKBL[88] NET_TRKBL[87] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_89 BL_TK VXDDAI VDDI VSSI WL[178] WL[179] TIEL FLOAT1[89] NET[89]
+ NET[88] NET_TRKBL[89] NET_TRKBL[88] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_90 BL_TK VXDDAI VDDI VSSI WL[180] WL[181] TIEL FLOAT1[90] NET[90]
+ NET[89] NET_TRKBL[90] NET_TRKBL[89] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_91 BL_TK VXDDAI VDDI VSSI WL[182] WL[183] TIEL FLOAT1[91] NET[91]
+ NET[90] NET_TRKBL[91] NET_TRKBL[90] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_92 BL_TK VXDDAI VDDI VSSI WL[184] WL[185] TIEL FLOAT1[92] NET[92]
+ NET[91] NET_TRKBL[92] NET_TRKBL[91] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_93 BL_TK VXDDAI VDDI VSSI WL[186] WL[187] TIEL FLOAT1[93] NET[93]
+ NET[92] NET_TRKBL[93] NET_TRKBL[92] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_94 BL_TK VXDDAI VDDI VSSI WL[188] WL[189] TIEL FLOAT1[94] NET[94]
+ NET[93] NET_TRKBL[94] NET_TRKBL[93] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_95 BL_TK VXDDAI VDDI VSSI WL[190] WL[191] TIEL FLOAT1[95] NET[95]
+ NET[94] NET_TRKBL[95] NET_TRKBL[94] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_96 BL_TK VXDDAI VDDI VSSI WL[192] WL[193] TIEL FLOAT1[96] NET[96]
+ NET[95] NET_TRKBL[96] NET_TRKBL[95] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_97 BL_TK VXDDAI VDDI VSSI WL[194] WL[195] TIEL FLOAT1[97] NET[97]
+ NET[96] NET_TRKBL[97] NET_TRKBL[96] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_98 BL_TK VXDDAI VDDI VSSI WL[196] WL[197] TIEL FLOAT1[98] NET[98]
+ NET[97] NET_TRKBL[98] NET_TRKBL[97] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_99 BL_TK VXDDAI VDDI VSSI WL[198] WL[199] TIEL FLOAT1[99] NET[99]
+ NET[98] NET_TRKBL[99] NET_TRKBL[98] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_100 BL_TK VXDDAI VDDI VSSI WL[200] WL[201] TIEL FLOAT1[100] NET[100]
+ NET[99] NET_TRKBL[100] NET_TRKBL[99] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_101 BL_TK VXDDAI VDDI VSSI WL[202] WL[203] TIEL FLOAT1[101] NET[101]
+ NET[100] NET_TRKBL[101] NET_TRKBL[100] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_102 BL_TK VXDDAI VDDI VSSI WL[204] WL[205] TIEL FLOAT1[102] NET[102]
+ NET[101] NET_TRKBL[102] NET_TRKBL[101] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_103 BL_TK VXDDAI VDDI VSSI WL[206] WL[207] TIEL FLOAT1[103] NET[103]
+ NET[102] NET_TRKBL[103] NET_TRKBL[102] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_104 BL_TK VXDDAI VDDI VSSI WL[208] WL[209] TIEL FLOAT1[104] NET[104]
+ NET[103] NET_TRKBL[104] NET_TRKBL[103] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_105 BL_TK VXDDAI VDDI VSSI WL[210] WL[211] TIEL FLOAT1[105] NET[105]
+ NET[104] NET_TRKBL[105] NET_TRKBL[104] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_106 BL_TK VXDDAI VDDI VSSI WL[212] WL[213] TIEL FLOAT1[106] NET[106]
+ NET[105] NET_TRKBL[106] NET_TRKBL[105] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_107 BL_TK VXDDAI VDDI VSSI WL[214] WL[215] TIEL FLOAT1[107] NET[107]
+ NET[106] NET_TRKBL[107] NET_TRKBL[106] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_108 BL_TK VXDDAI VDDI VSSI WL[216] WL[217] TIEL FLOAT1[108] NET[108]
+ NET[107] NET_TRKBL[108] NET_TRKBL[107] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_109 BL_TK VXDDAI VDDI VSSI WL[218] WL[219] TIEL FLOAT1[109] NET[109]
+ NET[108] NET_TRKBL[109] NET_TRKBL[108] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_110 BL_TK VXDDAI VDDI VSSI WL[220] WL[221] TIEL FLOAT1[110] NET[110]
+ NET[109] NET_TRKBL[110] NET_TRKBL[109] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_111 BL_TK VXDDAI VDDI VSSI WL[222] WL[223] TIEL FLOAT1[111] NET[111]
+ NET[110] NET_TRKBL[111] NET_TRKBL[110] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_112 BL_TK VXDDAI VDDI VSSI WL[224] WL[225] TIEL FLOAT1[112] NET[112]
+ NET[111] NET_TRKBL[112] NET_TRKBL[111] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_113 BL_TK VXDDAI VDDI VSSI WL[226] WL[227] TIEL FLOAT1[113] NET[113]
+ NET[112] NET_TRKBL[113] NET_TRKBL[112] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_114 BL_TK VXDDAI VDDI VSSI WL[228] WL[229] TIEL FLOAT1[114] NET[114]
+ NET[113] NET_TRKBL[114] NET_TRKBL[113] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_115 BL_TK VXDDAI VDDI VSSI WL[230] WL[231] TIEL FLOAT1[115] NET[115]
+ NET[114] NET_TRKBL[115] NET_TRKBL[114] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_116 BL_TK VXDDAI VDDI VSSI WL[232] WL[233] TIEL FLOAT1[116] NET[116]
+ NET[115] NET_TRKBL[116] NET_TRKBL[115] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_117 BL_TK VXDDAI VDDI VSSI WL[234] WL[235] TIEL FLOAT1[117] NET[117]
+ NET[116] NET_TRKBL[117] NET_TRKBL[116] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_118 BL_TK VXDDAI VDDI VSSI WL[236] WL[237] TIEL FLOAT1[118] NET[118]
+ NET[117] NET_TRKBL[118] NET_TRKBL[117] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_119 BL_TK VXDDAI VDDI VSSI WL[238] WL[239] TIEL FLOAT1[119] NET[119]
+ NET[118] NET_TRKBL[119] NET_TRKBL[118] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_120 BL_TK VXDDAI VDDI VSSI WL[240] WL[241] TIEL FLOAT1[120] NET[120]
+ NET[119] NET_TRKBL[120] NET_TRKBL[119] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_121 BL_TK VXDDAI VDDI VSSI WL[242] WL[243] TIEL FLOAT1[121] NET[121]
+ NET[120] NET_TRKBL[121] NET_TRKBL[120] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_122 BL_TK VXDDAI VDDI VSSI WL[244] WL[245] TIEL FLOAT1[122] NET[122]
+ NET[121] NET_TRKBL[122] NET_TRKBL[121] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_123 BL_TK VXDDAI VDDI VSSI WL[246] WL[247] TIEL FLOAT1[123] NET[123]
+ NET[122] NET_TRKBL[123] NET_TRKBL[122] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_124 BL_TK VXDDAI VDDI VSSI WL[248] WL[249] TIEL FLOAT1[124] NET[124]
+ NET[123] NET_TRKBL[124] NET_TRKBL[123] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_125 BL_TK VXDDAI VDDI VSSI WL[250] WL[251] TIEL FLOAT1[125] NET[125]
+ NET[124] NET_TRKBL[125] NET_TRKBL[124] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X4TRKNORX2_126 BL_TK VXDDAI VDDI VSSI WL[252] WL[253] TIEL FLOAT1[126] NET[126]
+ NET[125] NET_TRKBL[126] NET_TRKBL[125] TIEH S1BSVTSWSO8000Y24_TRKNORX2
X5TRKNORX2_127 BL_TK VXDDAI VDDI VSSI WL[254] WL[255] TIEL FLOAT1[127] NET[127]
+ NET[126] NET_TRKBL[127] NET_TRKBL[126] TIEH S1BSVTSWSO8000Y24_TRKNORX2
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_BANK_0_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6]
+ GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15]
+ GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23]
+ GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31]
+ GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6]
+ GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17]
+ GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28]
+ GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3]
+ GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13]
+ GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22]
+ GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31]
+ GWB[32] GWB[33] GWB[34] GWB[35] DSLP_BUF SLP_LCTRL RE WE VXDDHD WLP_SAE
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5]
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1]
+ DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] YL[1] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] BL_TK
+ WL_TK VXDDAI VDDI VSSI WLP_SAE_TK TK
XTRACKING WL_TK SLP_LCTRL BL_TK VXDDHD WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6]
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17]
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28]
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39]
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50]
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61]
+ WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72]
+ WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83]
+ WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94]
+ WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104]
+ WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113]
+ WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122]
+ WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] WL[131]
+ WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140]
+ WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149]
+ WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158]
+ WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167]
+ WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176]
+ WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185]
+ WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] WL[194]
+ WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203]
+ WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212]
+ WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221]
+ WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230]
+ WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239]
+ WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248]
+ WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] VXDDAI VDDI VSSI
+ S1BSVTSWSO8000Y24_TRACKING
XLIO_MCB_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] VXDDAI LIOPD WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7]
+ WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18]
+ WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29]
+ WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40]
+ WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51]
+ WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62]
+ WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73]
+ WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84]
+ WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95]
+ WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105]
+ WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114]
+ WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123]
+ WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] WL[132]
+ WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141]
+ WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150]
+ WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159]
+ WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168]
+ WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177]
+ WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186]
+ WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] WL[195]
+ WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204]
+ WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213]
+ WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222]
+ WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231]
+ WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240]
+ WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249]
+ WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] WL[258]
+ WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] WL[267]
+ WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] WL[276]
+ WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] WL[285]
+ WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] WL[294]
+ WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] WL[303]
+ WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] WL[312]
+ WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] WL[321]
+ WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] WL[330]
+ WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] WL[339]
+ WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] WL[348]
+ WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] WL[357]
+ WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] WL[366]
+ WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] WL[375]
+ WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] WL[383] WL[384]
+ WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] WL[392] WL[393]
+ WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] WL[401] WL[402]
+ WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] WL[410] WL[411]
+ WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] WL[419] WL[420]
+ WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] WL[428] WL[429]
+ WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] WL[437] WL[438]
+ WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] WL[446] WL[447]
+ WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] WL[455] WL[456]
+ WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] WL[464] WL[465]
+ WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] WL[473] WL[474]
+ WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] WL[482] WL[483]
+ WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] WL[491] WL[492]
+ WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] WL[500] WL[501]
+ WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] WL[509] WL[510]
+ WL[511] BLEQ_DN BLEQ_UP GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8]
+ GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19]
+ GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30]
+ GW[31] GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5]
+ GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15]
+ GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24]
+ GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33]
+ GWB[34] GWB[35] RE_LIO SAEB WE_LIO DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2]
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0]
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6]
+ DEC_Y_UP[7] YL_LIO[0] YL_LIO[1] VDDI VSSI S1BSVTSWSO8000Y24_LIO_MCB_F
XLCTRL_S_M16_SD BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1]
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4]
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4]
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3]
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1]
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7]
+ DSLP_BUF LIOPD RE RE_LIO SAEB SLP_LCTRL TK VXDDHD VDDI VSSI WE WE_LIO
+ WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2]
+ WLPY_UP[3] WLP_SAE WLP_SAE_TK YL[0] YL[1] YL_LIO[0] YL_LIO[1]
+ S1BSVTSWSO8000Y24_LCTRL_S_M16_SD
XXDRV_STRAPD0 VXDDHD VDDI VSSI WLPY_DN[0] WLPY_DNB[0]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_SHA_0 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD0 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[0] WL[1]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_1 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD0 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[2] WL[3]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS1 DEC_X1[0] SH_NPD0 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_2 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD1 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[4] WL[5]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_3 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD1 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[6] WL[7]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS3 DEC_X1[0] SH_NPD1 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_4 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD2 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[8] WL[9]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_5 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD2 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[10] WL[11]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS5 DEC_X1[1] SH_NPD2 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_6 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD3 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[12] WL[13]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_7 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD3 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[14] WL[15]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS7 DEC_X1[1] SH_NPD3 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_8 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD4 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[16] WL[17]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_9 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD4 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[18] WL[19]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS9 DEC_X1[2] SH_NPD4 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_10 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD5 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[20] WL[21]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_11 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD5 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[22] WL[23]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS11 DEC_X1[2] SH_NPD5 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_12 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD6 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[24] WL[25]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_13 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD6 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[26] WL[27]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS13 DEC_X1[3] SH_NPD6 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_14 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD7 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[28] WL[29]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_15 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD7 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[30] WL[31]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS15 DEC_X1[3] SH_NPD7 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_16 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD8 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[32] WL[33]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_17 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD8 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[34] WL[35]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS17 DEC_X1[4] SH_NPD8 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_18 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD9 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[36] WL[37]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_19 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD9 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[38] WL[39]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS19 DEC_X1[4] SH_NPD9 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_20 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD10 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[40] WL[41]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_21 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD10 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[42] WL[43]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS21 DEC_X1[5] SH_NPD10 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_22 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD11 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[44] WL[45]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_23 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD11 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[46] WL[47]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS23 DEC_X1[5] SH_NPD11 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_24 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD12 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[48] WL[49]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_25 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD12 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[50] WL[51]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS25 DEC_X1[6] SH_NPD12 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_26 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD13 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[52] WL[53]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_27 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD13 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[54] WL[55]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS27 DEC_X1[6] SH_NPD13 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_28 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD14 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[56] WL[57]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_29 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD14 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[58] WL[59]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS29 DEC_X1[7] SH_NPD14 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_30 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD15 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[60] WL[61]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_31 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD15 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[62] WL[63]
+ WLPY_DN[0] WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS31 DEC_X1[7] SH_NPD15 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPD1 VXDDHD VDDI VSSI WLPY_DN[1] WLPY_DNB[1]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_SHA_32 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD16 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[64] WL[65]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_33 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD16 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[66] WL[67]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS33 DEC_X1[0] SH_NPD16 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_34 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD17 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[68] WL[69]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_35 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD17 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[70] WL[71]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS35 DEC_X1[0] SH_NPD17 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_36 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD18 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[72] WL[73]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_37 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD18 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[74] WL[75]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS37 DEC_X1[1] SH_NPD18 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_38 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD19 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[76] WL[77]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_39 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD19 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[78] WL[79]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS39 DEC_X1[1] SH_NPD19 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_40 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD20 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[80] WL[81]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_41 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD20 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[82] WL[83]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS41 DEC_X1[2] SH_NPD20 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_42 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD21 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[84] WL[85]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_43 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD21 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[86] WL[87]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS43 DEC_X1[2] SH_NPD21 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_44 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD22 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[88] WL[89]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_45 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD22 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[90] WL[91]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS45 DEC_X1[3] SH_NPD22 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_46 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD23 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[92] WL[93]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_47 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD23 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[94] WL[95]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS47 DEC_X1[3] SH_NPD23 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_48 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD24 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[96] WL[97]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_49 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD24 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[98] WL[99]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS49 DEC_X1[4] SH_NPD24 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_50 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD25 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[100] WL[101]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_51 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD25 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[102] WL[103]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS51 DEC_X1[4] SH_NPD25 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_52 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD26 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[104] WL[105]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_53 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD26 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[106] WL[107]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS53 DEC_X1[5] SH_NPD26 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_54 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD27 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[108] WL[109]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_55 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD27 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[110] WL[111]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS55 DEC_X1[5] SH_NPD27 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_56 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD28 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[112] WL[113]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_57 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD28 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[114] WL[115]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS57 DEC_X1[6] SH_NPD28 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_58 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD29 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[116] WL[117]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_59 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD29 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[118] WL[119]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS59 DEC_X1[6] SH_NPD29 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_60 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD30 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[120] WL[121]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_61 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD30 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[122] WL[123]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS61 DEC_X1[7] SH_NPD30 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_62 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD31 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[124] WL[125]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_63 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD31 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[126] WL[127]
+ WLPY_DN[1] WLPY_DNB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS63 DEC_X1[7] SH_NPD31 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPD2 VXDDHD VDDI VSSI WLPY_DN[2] WLPY_DNB[2]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_SHA_64 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD32 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[128] WL[129]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_65 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD32 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[130] WL[131]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS65 DEC_X1[0] SH_NPD32 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_66 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD33 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[132] WL[133]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_67 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD33 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[134] WL[135]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS67 DEC_X1[0] SH_NPD33 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_68 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD34 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[136] WL[137]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_69 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD34 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[138] WL[139]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS69 DEC_X1[1] SH_NPD34 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_70 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD35 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[140] WL[141]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_71 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD35 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[142] WL[143]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS71 DEC_X1[1] SH_NPD35 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_72 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD36 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[144] WL[145]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_73 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD36 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[146] WL[147]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS73 DEC_X1[2] SH_NPD36 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_74 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD37 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[148] WL[149]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_75 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD37 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[150] WL[151]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS75 DEC_X1[2] SH_NPD37 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_76 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD38 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[152] WL[153]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_77 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD38 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[154] WL[155]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS77 DEC_X1[3] SH_NPD38 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_78 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD39 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[156] WL[157]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_79 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD39 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[158] WL[159]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS79 DEC_X1[3] SH_NPD39 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_80 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD40 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[160] WL[161]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_81 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD40 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[162] WL[163]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS81 DEC_X1[4] SH_NPD40 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_82 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD41 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[164] WL[165]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_83 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD41 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[166] WL[167]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS83 DEC_X1[4] SH_NPD41 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_84 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD42 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[168] WL[169]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_85 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD42 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[170] WL[171]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS85 DEC_X1[5] SH_NPD42 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_86 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD43 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[172] WL[173]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_87 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD43 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[174] WL[175]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS87 DEC_X1[5] SH_NPD43 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_88 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD44 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[176] WL[177]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_89 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD44 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[178] WL[179]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS89 DEC_X1[6] SH_NPD44 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_90 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD45 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[180] WL[181]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_91 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD45 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[182] WL[183]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS91 DEC_X1[6] SH_NPD45 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_92 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD46 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[184] WL[185]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_93 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD46 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[186] WL[187]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS93 DEC_X1[7] SH_NPD46 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_94 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD47 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[188] WL[189]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_95 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD47 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[190] WL[191]
+ WLPY_DN[2] WLPY_DNB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS95 DEC_X1[7] SH_NPD47 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPD3 VXDDHD VDDI VSSI WLPY_DN[3] WLPY_DNB[3]
+ S1BSVTSWSO8000Y24_XDRV_STRAP_LCNT
XXDRV_LA512_SHA_96 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD48 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[192] WL[193]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_97 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD48 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[194] WL[195]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS97 DEC_X1[0] SH_NPD48 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_98 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD49 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[196] WL[197]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_99 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD49 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[198] WL[199]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS99 DEC_X1[0] SH_NPD49 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_100 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD50 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[200] WL[201]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_101 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD50 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[202] WL[203]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS101 DEC_X1[1] SH_NPD50 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_102 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD51 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[204] WL[205]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_103 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD51 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[206] WL[207]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS103 DEC_X1[1] SH_NPD51 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_104 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD52 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[208] WL[209]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_105 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD52 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[210] WL[211]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS105 DEC_X1[2] SH_NPD52 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_106 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD53 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[212] WL[213]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_107 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD53 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[214] WL[215]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS107 DEC_X1[2] SH_NPD53 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_108 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD54 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[216] WL[217]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_109 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD54 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[218] WL[219]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS109 DEC_X1[3] SH_NPD54 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_110 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD55 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[220] WL[221]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_111 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD55 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[222] WL[223]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS111 DEC_X1[3] SH_NPD55 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_112 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD56 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[224] WL[225]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_113 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD56 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[226] WL[227]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS113 DEC_X1[4] SH_NPD56 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_114 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD57 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[228] WL[229]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_115 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD57 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[230] WL[231]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS115 DEC_X1[4] SH_NPD57 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_116 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD58 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[232] WL[233]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_117 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD58 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[234] WL[235]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS117 DEC_X1[5] SH_NPD58 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_118 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD59 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[236] WL[237]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_119 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD59 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[238] WL[239]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS119 DEC_X1[5] SH_NPD59 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_120 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD60 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[240] WL[241]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_121 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD60 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[242] WL[243]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS121 DEC_X1[6] SH_NPD60 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_122 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD61 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[244] WL[245]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_123 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD61 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[246] WL[247]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS123 DEC_X1[6] SH_NPD61 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_124 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD62 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[248] WL[249]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_125 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD62 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[250] WL[251]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS125 DEC_X1[7] SH_NPD62 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_126 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD63 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[252] WL[253]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_127 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD63 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[254] WL[255]
+ WLPY_DN[3] WLPY_DNB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS127 DEC_X1[7] SH_NPD63 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPU0 VXDDHD VDDI VSSI WLPY_UP[0] WLPY_UPB[0]
+ S1BSVTSWSO8000Y24_XDRV_STRAP_LCNT
XXDRV_LA512_SHA_128 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD64 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[256] WL[257]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_129 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD64 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[258] WL[259]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS129 DEC_X1[0] SH_NPD64 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_130 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD65 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[260] WL[261]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_131 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD65 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[262] WL[263]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS131 DEC_X1[0] SH_NPD65 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_132 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD66 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[264] WL[265]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_133 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD66 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[266] WL[267]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS133 DEC_X1[1] SH_NPD66 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_134 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD67 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[268] WL[269]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_135 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD67 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[270] WL[271]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS135 DEC_X1[1] SH_NPD67 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_136 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD68 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[272] WL[273]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_137 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD68 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[274] WL[275]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS137 DEC_X1[2] SH_NPD68 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_138 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD69 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[276] WL[277]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_139 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD69 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[278] WL[279]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS139 DEC_X1[2] SH_NPD69 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_140 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD70 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[280] WL[281]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_141 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD70 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[282] WL[283]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS141 DEC_X1[3] SH_NPD70 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_142 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD71 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[284] WL[285]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_143 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD71 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[286] WL[287]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS143 DEC_X1[3] SH_NPD71 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_144 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD72 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[288] WL[289]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_145 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD72 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[290] WL[291]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS145 DEC_X1[4] SH_NPD72 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_146 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD73 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[292] WL[293]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_147 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD73 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[294] WL[295]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS147 DEC_X1[4] SH_NPD73 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_148 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD74 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[296] WL[297]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_149 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD74 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[298] WL[299]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS149 DEC_X1[5] SH_NPD74 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_150 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD75 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[300] WL[301]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_151 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD75 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[302] WL[303]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS151 DEC_X1[5] SH_NPD75 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_152 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD76 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[304] WL[305]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_153 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD76 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[306] WL[307]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS153 DEC_X1[6] SH_NPD76 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_154 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD77 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[308] WL[309]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_155 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD77 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[310] WL[311]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS155 DEC_X1[6] SH_NPD77 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_156 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD78 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[312] WL[313]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_157 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD78 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[314] WL[315]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS157 DEC_X1[7] SH_NPD78 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_158 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD79 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[316] WL[317]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_159 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD79 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[318] WL[319]
+ WLPY_UP[0] WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS159 DEC_X1[7] SH_NPD79 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPU1 VXDDHD VDDI VSSI WLPY_UP[1] WLPY_UPB[1]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_SHA_160 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD80 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[320] WL[321]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_161 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD80 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[322] WL[323]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS161 DEC_X1[0] SH_NPD80 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_162 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD81 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[324] WL[325]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_163 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD81 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[326] WL[327]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS163 DEC_X1[0] SH_NPD81 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_164 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD82 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[328] WL[329]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_165 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD82 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[330] WL[331]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS165 DEC_X1[1] SH_NPD82 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_166 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD83 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[332] WL[333]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_167 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD83 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[334] WL[335]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS167 DEC_X1[1] SH_NPD83 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_168 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD84 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[336] WL[337]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_169 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD84 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[338] WL[339]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS169 DEC_X1[2] SH_NPD84 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_170 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD85 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[340] WL[341]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_171 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD85 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[342] WL[343]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS171 DEC_X1[2] SH_NPD85 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_172 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD86 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[344] WL[345]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_173 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD86 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[346] WL[347]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS173 DEC_X1[3] SH_NPD86 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_174 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD87 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[348] WL[349]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_175 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD87 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[350] WL[351]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS175 DEC_X1[3] SH_NPD87 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_176 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD88 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[352] WL[353]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_177 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD88 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[354] WL[355]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS177 DEC_X1[4] SH_NPD88 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_178 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD89 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[356] WL[357]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_179 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD89 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[358] WL[359]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS179 DEC_X1[4] SH_NPD89 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_180 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD90 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[360] WL[361]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_181 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD90 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[362] WL[363]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS181 DEC_X1[5] SH_NPD90 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_182 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD91 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[364] WL[365]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_183 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD91 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[366] WL[367]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS183 DEC_X1[5] SH_NPD91 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_184 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD92 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[368] WL[369]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_185 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD92 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[370] WL[371]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS185 DEC_X1[6] SH_NPD92 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_186 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD93 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[372] WL[373]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_187 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD93 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[374] WL[375]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS187 DEC_X1[6] SH_NPD93 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_188 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD94 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[376] WL[377]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_189 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD94 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[378] WL[379]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS189 DEC_X1[7] SH_NPD94 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_190 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD95 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[380] WL[381]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_191 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD95 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[382] WL[383]
+ WLPY_UP[1] WLPY_UPB[1] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS191 DEC_X1[7] SH_NPD95 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPU2 VXDDHD VDDI VSSI WLPY_UP[2] WLPY_UPB[2]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_SHA_192 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD96 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[384] WL[385]
+ WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_193 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD96 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[386] WL[387]
+ WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS193 DEC_X1[0] SH_NPD96 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_194 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD97 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[388] WL[389]
+ WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_195 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD97 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[390] WL[391]
+ WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS195 DEC_X1[0] SH_NPD97 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_196 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD98 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[392] WL[393]
+ WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_197 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD98 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[394] WL[395]
+ WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS197 DEC_X1[1] SH_NPD98 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_198 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD99 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[396] WL[397]
+ WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_199 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD99 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[398] WL[399]
+ WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS199 DEC_X1[1] SH_NPD99 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_200 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD100 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[400]
+ WL[401] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_201 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD100 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[402]
+ WL[403] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS201 DEC_X1[2] SH_NPD100 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_202 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD101 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[404]
+ WL[405] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_203 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD101 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[406]
+ WL[407] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS203 DEC_X1[2] SH_NPD101 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_204 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD102 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[408]
+ WL[409] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_205 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD102 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[410]
+ WL[411] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS205 DEC_X1[3] SH_NPD102 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_206 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD103 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[412]
+ WL[413] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_207 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD103 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[414]
+ WL[415] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS207 DEC_X1[3] SH_NPD103 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_208 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD104 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[416]
+ WL[417] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_209 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD104 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[418]
+ WL[419] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS209 DEC_X1[4] SH_NPD104 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_210 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD105 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[420]
+ WL[421] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_211 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD105 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[422]
+ WL[423] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS211 DEC_X1[4] SH_NPD105 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_212 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD106 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[424]
+ WL[425] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_213 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD106 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[426]
+ WL[427] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS213 DEC_X1[5] SH_NPD106 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_214 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD107 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[428]
+ WL[429] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_215 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD107 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[430]
+ WL[431] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS215 DEC_X1[5] SH_NPD107 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_216 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD108 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[432]
+ WL[433] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_217 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD108 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[434]
+ WL[435] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS217 DEC_X1[6] SH_NPD108 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_218 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD109 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[436]
+ WL[437] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_219 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD109 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[438]
+ WL[439] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS219 DEC_X1[6] SH_NPD109 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_220 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD110 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[440]
+ WL[441] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_221 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD110 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[442]
+ WL[443] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS221 DEC_X1[7] SH_NPD110 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_222 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD111 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[444]
+ WL[445] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_223 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD111 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[446]
+ WL[447] WLPY_UP[2] WLPY_UPB[2] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS223 DEC_X1[7] SH_NPD111 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_STRAPU3 VXDDHD VDDI VSSI WLPY_UP[3] WLPY_UPB[3]
+ S1BSVTSWSO8000Y24_XDRV_STRAP
XXDRV_LA512_SHA_224 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD112 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[448]
+ WL[449] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_225 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD112 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[450]
+ WL[451] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS225 DEC_X1[0] SH_NPD112 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_226 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD113 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[452]
+ WL[453] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_227 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD113 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[454]
+ WL[455] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS227 DEC_X1[0] SH_NPD113 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_228 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD114 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[456]
+ WL[457] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_229 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD114 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[458]
+ WL[459] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS229 DEC_X1[1] SH_NPD114 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_230 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD115 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[460]
+ WL[461] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_231 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD115 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[462]
+ WL[463] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS231 DEC_X1[1] SH_NPD115 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_232 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD116 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[464]
+ WL[465] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_233 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD116 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[466]
+ WL[467] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS233 DEC_X1[2] SH_NPD116 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_234 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD117 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[468]
+ WL[469] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_235 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD117 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[470]
+ WL[471] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS235 DEC_X1[2] SH_NPD117 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_236 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD118 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[472]
+ WL[473] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_237 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD118 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[474]
+ WL[475] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS237 DEC_X1[3] SH_NPD118 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_238 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD119 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[476]
+ WL[477] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_239 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD119 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[478]
+ WL[479] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS239 DEC_X1[3] SH_NPD119 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_240 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD120 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[480]
+ WL[481] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_241 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD120 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[482]
+ WL[483] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS241 DEC_X1[4] SH_NPD120 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_242 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD121 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[484]
+ WL[485] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_243 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD121 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[486]
+ WL[487] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS243 DEC_X1[4] SH_NPD121 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_244 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD122 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[488]
+ WL[489] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_245 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD122 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[490]
+ WL[491] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS245 DEC_X1[5] SH_NPD122 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_246 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD123 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[492]
+ WL[493] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_247 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD123 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[494]
+ WL[495] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS247 DEC_X1[5] SH_NPD123 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_248 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD124 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[496]
+ WL[497] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_249 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD124 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[498]
+ WL[499] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS249 DEC_X1[6] SH_NPD124 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_250 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD125 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[500]
+ WL[501] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_251 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD125 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[502]
+ WL[503] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS251 DEC_X1[6] SH_NPD125 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_252 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD126 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[504]
+ WL[505] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_253 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD126 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[506]
+ WL[507] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS253 DEC_X1[7] SH_NPD126 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
XXDRV_LA512_SHA_254 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD127 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[508]
+ WL[509] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_255 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] DSLP_BUF RE SH_NPD127 SLP_LCTRL TK VXDDHD VDDI VSSI WE WL[510]
+ WL[511] WLPY_UP[3] WLPY_UPB[3] WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA
XXDRV_LA512_SHA_NMOS255 DEC_X1[7] SH_NPD127 VSSI
+ S1BSVTSWSO8000Y24_XDRV_LA512_SHA_NMOS
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_CNT_CORE_IO_DR AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB
+ CEBM CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] RTSEL[0] RTSEL[1] RE WE TK TM TRKBL VXDDFHD VDDF VHI VLO VSSI WEB
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2]
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5]
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1]
+ YM[2] YM[3] DSLP DSLP_BUF SD SD_BUF SLP SLP_BUF SLP_LBACK SLP_LCTRL SLP_Q
+ SLP_RBACK BWEB[0] BWEB[1] BWEBM[0] BWEBM[1] D[0] D[1] DM[0] DM[1] GBL[0]
+ GBL[1] GBLB[0] GBLB[1] GW[0] GW[1] GWB[0] GWB[1] Q[0] Q[1] VXDDHD VDDI
+ SLP_VXDD VLO_VXDD VHI_VXDD
XCNT_M16_IOX2_WOBIST_SR AWT AWT2 BLTRKWLDRV BWEB[0] BWEB[1] CEB CKD CLK
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5]
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF D[0]
+ D[1] GBLB[0] GBLB[1] GBL[0] GBL[1] GWB[0] GWB[1] GW[0] GW[1] Q[0] Q[1] RE
+ RTSEL[0] RTSEL[1] SD SLP SLP_BUF SLP_LBACK SLP_LCTRL SLP_Q SLP_RBACK TK TM
+ TRKBL VXDDHD VDDI VHI VHI_VXDD VLO VLO_VXDD VSSI WE WEB WLP_SAE WLP_SAEB
+ WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7]
+ X[8] X[9] X[10] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1]
+ S1BSVTSWSO8000Y24_CNT_M16_IOX2_WOBIST_SR
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_MIO_L_DR AWT BIST BWEB[0] BWEB[1] BWEB[2] BWEB[3]
+ BWEB[4] BWEB[5] BWEB[6] BWEB[7] BWEB[8] BWEB[9] BWEB[10] BWEB[11] BWEB[12]
+ BWEB[13] BWEB[14] BWEB[15] BWEB[16] BWEBM[0] BWEBM[1] BWEBM[2] BWEBM[3]
+ BWEBM[4] BWEBM[5] BWEBM[6] BWEBM[7] BWEBM[8] BWEBM[9] BWEBM[10] BWEBM[11]
+ BWEBM[12] BWEBM[13] BWEBM[14] BWEBM[15] BWEBM[16] CKD D[0] D[1] D[2] D[3] D[4]
+ D[5] D[6] D[7] D[8] D[9] D[10] D[11] D[12] D[13] D[14] D[15] D[16] DM[0] DM[1]
+ DM[2] DM[3] DM[4] DM[5] DM[6] DM[7] DM[8] DM[9] DM[10] DM[11] DM[12] DM[13]
+ DM[14] DM[15] DM[16] GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7]
+ GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GW[0] GW[1]
+ GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13]
+ GW[14] GW[15] GW[16] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] IOPD PDI
+ PDO Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] Q[10] Q[11] Q[12] Q[13]
+ Q[14] Q[15] Q[16] SLP_Q VXDDHD VDDF VSSI VLO WLP_SAEB PDOL[2] CVXDDHD VDDI
+ SLP_VXDD VXDDFHD
XIO_M16_0 AWT BWEB[0] CKD D[0] GBL[0] GBLB[0] GW[0] GWB[0] IOPD PDI PDOL[0] Q[0]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16_WOBIST_SR
XIO_M16B_1 AWT BWEB[1] CKD D[1] GBL[1] GBLB[1] GW[1] GWB[1] PDOL[0] Q[1] SLP_Q
+ VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_2 AWT BWEB[2] CKD D[2] GBL[2] GBLB[2] GW[2] GWB[2] PDOL[0] Q[2] SLP_Q
+ VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_3 AWT BWEB[3] CKD D[3] GBL[3] GBLB[3] GW[3] GWB[3] PDOL[0] Q[3] SLP_Q
+ VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_4 AWT BWEB[4] CKD D[4] GBL[4] GBLB[4] GW[4] GWB[4] PDOL[0] Q[4] SLP_Q
+ VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_5 AWT BWEB[5] CKD D[5] GBL[5] GBLB[5] GW[5] GWB[5] PDOL[0] Q[5] SLP_Q
+ VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_6 AWT BWEB[6] CKD D[6] GBL[6] GBLB[6] GW[6] GWB[6] PDOL[0] Q[6] SLP_Q
+ VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_7 AWT BWEB[7] CKD D[7] GBL[7] GBLB[7] GW[7] GWB[7] PDOL[0] Q[7] SLP_Q
+ VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16_8 AWT BWEB[8] CKD D[8] GBL[8] GBLB[8] GW[8] GWB[8] IOPD PDOL[0] PDOL[1]
+ Q[8] SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16_WOBIST_SR
XIO_M16B_9 AWT BWEB[9] CKD D[9] GBL[9] GBLB[9] GW[9] GWB[9] PDOL[1] Q[9] SLP_Q
+ VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_10 AWT BWEB[10] CKD D[10] GBL[10] GBLB[10] GW[10] GWB[10] PDOL[1] Q[10]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_11 AWT BWEB[11] CKD D[11] GBL[11] GBLB[11] GW[11] GWB[11] PDOL[1] Q[11]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_12 AWT BWEB[12] CKD D[12] GBL[12] GBLB[12] GW[12] GWB[12] PDOL[1] Q[12]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_13 AWT BWEB[13] CKD D[13] GBL[13] GBLB[13] GW[13] GWB[13] PDOL[1] Q[13]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_14 AWT BWEB[14] CKD D[14] GBL[14] GBLB[14] GW[14] GWB[14] PDOL[1] Q[14]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_15 AWT BWEB[15] CKD D[15] GBL[15] GBLB[15] GW[15] GWB[15] PDOL[1] Q[15]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16_16 AWT BWEB[16] CKD D[16] GBL[16] GBLB[16] GW[16] GWB[16] IOPD PDOL[1]
+ PDOL[2] Q[16] SLP_Q VXDDHD VDDI VSSI WLP_SAEB
+ S1BSVTSWSO8000Y24_IO_M16_WOBIST_SR
.ENDS

.SUBCKT S1BSVTSWSO8000Y24_MIO_R_DR AWT BIST BWEB[19] BWEB[20] BWEB[21] BWEB[22]
+ BWEB[23] BWEB[24] BWEB[25] BWEB[26] BWEB[27] BWEB[28] BWEB[29] BWEB[30]
+ BWEB[31] BWEB[32] BWEB[33] BWEB[34] BWEB[35] BWEBM[19] BWEBM[20] BWEBM[21]
+ BWEBM[22] BWEBM[23] BWEBM[24] BWEBM[25] BWEBM[26] BWEBM[27] BWEBM[28]
+ BWEBM[29] BWEBM[30] BWEBM[31] BWEBM[32] BWEBM[33] BWEBM[34] BWEBM[35] CKD
+ D[19] D[20] D[21] D[22] D[23] D[24] D[25] D[26] D[27] D[28] D[29] D[30] D[31]
+ D[32] D[33] D[34] D[35] DM[19] DM[20] DM[21] DM[22] DM[23] DM[24] DM[25]
+ DM[26] DM[27] DM[28] DM[29] DM[30] DM[31] DM[32] DM[33] DM[34] DM[35] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[19] GBLB[20]
+ GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28]
+ GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[19] GW[20]
+ GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31]
+ GW[32] GW[33] GW[34] GW[35] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24]
+ GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33]
+ GWB[34] GWB[35] IOPD PDI PDO Q[19] Q[20] Q[21] Q[22] Q[23] Q[24] Q[25] Q[26]
+ Q[27] Q[28] Q[29] Q[30] Q[31] Q[32] Q[33] Q[34] Q[35] SLP_Q VXDDHD VDDF VSSI
+ VLO WLP_SAEB PDOR[2] CVXDDHD VDDI SLP_VXDD VXDDFHD
XIO_M16_19 AWT BWEB[19] CKD D[19] GBL[19] GBLB[19] GW[19] GWB[19] IOPD PDI
+ PDOR[0] Q[19] SLP_Q VXDDHD VDDI VSSI WLP_SAEB
+ S1BSVTSWSO8000Y24_IO_M16_WOBIST_SR
XIO_M16B_20 AWT BWEB[20] CKD D[20] GBL[20] GBLB[20] GW[20] GWB[20] PDOR[0] Q[20]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_21 AWT BWEB[21] CKD D[21] GBL[21] GBLB[21] GW[21] GWB[21] PDOR[0] Q[21]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_22 AWT BWEB[22] CKD D[22] GBL[22] GBLB[22] GW[22] GWB[22] PDOR[0] Q[22]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_23 AWT BWEB[23] CKD D[23] GBL[23] GBLB[23] GW[23] GWB[23] PDOR[0] Q[23]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_24 AWT BWEB[24] CKD D[24] GBL[24] GBLB[24] GW[24] GWB[24] PDOR[0] Q[24]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_25 AWT BWEB[25] CKD D[25] GBL[25] GBLB[25] GW[25] GWB[25] PDOR[0] Q[25]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_26 AWT BWEB[26] CKD D[26] GBL[26] GBLB[26] GW[26] GWB[26] PDOR[0] Q[26]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16_27 AWT BWEB[27] CKD D[27] GBL[27] GBLB[27] GW[27] GWB[27] IOPD PDOR[0]
+ PDOR[1] Q[27] SLP_Q VXDDHD VDDI VSSI WLP_SAEB
+ S1BSVTSWSO8000Y24_IO_M16_WOBIST_SR
XIO_M16B_28 AWT BWEB[28] CKD D[28] GBL[28] GBLB[28] GW[28] GWB[28] PDOR[1] Q[28]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_29 AWT BWEB[29] CKD D[29] GBL[29] GBLB[29] GW[29] GWB[29] PDOR[1] Q[29]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_30 AWT BWEB[30] CKD D[30] GBL[30] GBLB[30] GW[30] GWB[30] PDOR[1] Q[30]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_31 AWT BWEB[31] CKD D[31] GBL[31] GBLB[31] GW[31] GWB[31] PDOR[1] Q[31]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_32 AWT BWEB[32] CKD D[32] GBL[32] GBLB[32] GW[32] GWB[32] PDOR[1] Q[32]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_33 AWT BWEB[33] CKD D[33] GBL[33] GBLB[33] GW[33] GWB[33] PDOR[1] Q[33]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16B_34 AWT BWEB[34] CKD D[34] GBL[34] GBLB[34] GW[34] GWB[34] PDOR[1] Q[34]
+ SLP_Q VXDDHD VDDI VSSI WLP_SAEB S1BSVTSWSO8000Y24_IO_M16B_WOBIST_SR
XIO_M16_35 AWT BWEB[35] CKD D[35] GBL[35] GBLB[35] GW[35] GWB[35] IOPD PDOR[1]
+ PDOR[2] Q[35] SLP_Q VXDDHD VDDI VSSI WLP_SAEB
+ S1BSVTSWSO8000Y24_IO_M16_WOBIST_SR
.ENDS

.SUBCKT TS1N28HPCPSVTB32768X36M16SWSO Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7]
+ Q[8] Q[9] Q[10] Q[11] Q[12] Q[13] Q[14] Q[15] Q[16] Q[17] Q[18] Q[19] Q[20]
+ Q[21] Q[22] Q[23] Q[24] Q[25] Q[26] Q[27] Q[28] Q[29] Q[30] Q[31] Q[32] Q[33]
+ Q[34] Q[35] A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] A[8] A[9] A[10] A[11]
+ A[12] A[13] A[14] BWEB[0] BWEB[1] BWEB[2] BWEB[3] BWEB[4] BWEB[5] BWEB[6]
+ BWEB[7] BWEB[8] BWEB[9] BWEB[10] BWEB[11] BWEB[12] BWEB[13] BWEB[14] BWEB[15]
+ BWEB[16] BWEB[17] BWEB[18] BWEB[19] BWEB[20] BWEB[21] BWEB[22] BWEB[23]
+ BWEB[24] BWEB[25] BWEB[26] BWEB[27] BWEB[28] BWEB[29] BWEB[30] BWEB[31]
+ BWEB[32] BWEB[33] BWEB[34] BWEB[35] CEB CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6]
+ D[7] D[8] D[9] D[10] D[11] D[12] D[13] D[14] D[15] D[16] D[17] D[18] D[19]
+ D[20] D[21] D[22] D[23] D[24] D[25] D[26] D[27] D[28] D[29] D[30] D[31] D[32]
+ D[33] D[34] D[35] SLP SD WEB VDD VSS
XBANK_0 GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9]
+ GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20]
+ GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31]
+ GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] DSLP_BUF SLP_LCTRL RE WE VXDDHD WLP_SAE DEC_X0[0] DEC_X0[1] DEC_X0[2]
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1]
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0]
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4]
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] YL[1] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3]
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] TRKBL BLTRKWLDRV VXDDAI VDD VSS
+ WLP_SAE_TK TK S1BSVTSWSO8000Y24_BANK_0_F
XREPEATER DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3]
+ DEC_X0_REP[4] DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1[0] DEC_X1[1]
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X1_REP[0]
+ DEC_X1_REP[1] DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5]
+ DEC_X1_REP[6] DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DSLP_BUF RE
+ SLP_LCTRL SLP_LCTRL_REP TK VXDDHD VDD VSS WE WLP_SAE WLP_SAE_TK YL[0] YL[1]
+ S1BSVTSWSO8000Y24_REPEATER
XBANK_1 GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9]
+ GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20]
+ GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31]
+ GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] DSLP_BUF SLP_LCTRL SLP_LCTRL_REP RE WE VXDDHD WLP_SAE DEC_X0[0]
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7]
+ DEC_X0_REP[0] DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4]
+ DEC_X0_REP[5] DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1[0] DEC_X1[1] DEC_X1[2]
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X1_REP[0] DEC_X1_REP[1]
+ DEC_X1_REP[2] DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5] DEC_X1_REP[6]
+ DEC_X1_REP[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1]
+ DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] YL[1] DEC_X3[2]
+ DEC_X3[3] DEC_X3[0] DEC_X3[1] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] VXDDAI
+ VDD VSS WLP_SAE_TK TK S1BSVTSWSO8000Y24_BANK_F_UP_REP
XBANK_2 GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9]
+ GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20]
+ GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31]
+ GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] DSLP_BUF SLP_LCTRL_REP RE WE VXDDHD WLP_SAE DEC_X0_REP[0]
+ DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5]
+ DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2]
+ DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5] DEC_X1_REP[6] DEC_X1_REP[7]
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3]
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] YL[1] DEC_X3[4] DEC_X3[5] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[6] DEC_X3[7] VXDDAI VDD VSS WLP_SAE_TK TK
+ S1BSVTSWSO8000Y24_BANK_F_REP
XBANK_3 GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9]
+ GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20]
+ GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31]
+ GW[32] GW[33] GW[34] GW[35] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] DSLP_BUF SLP_LCTRL_REP RE WE VXDDHD WLP_SAE DEC_X0_REP[0]
+ DEC_X0_REP[1] DEC_X0_REP[2] DEC_X0_REP[3] DEC_X0_REP[4] DEC_X0_REP[5]
+ DEC_X0_REP[6] DEC_X0_REP[7] DEC_X1_REP[0] DEC_X1_REP[1] DEC_X1_REP[2]
+ DEC_X1_REP[3] DEC_X1_REP[4] DEC_X1_REP[5] DEC_X1_REP[6] DEC_X1_REP[7]
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3]
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] YL[1] DEC_X3[6] DEC_X3[7] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] VXDDAI VDD VSS WLP_SAE_TK TK
+ S1BSVTSWSO8000Y24_BANK_F_REP
XMIO_L AWT2 VLO_VXDD BWEB[0] BWEB[1] BWEB[2] BWEB[3] BWEB[4] BWEB[5] BWEB[6]
+ BWEB[7] BWEB[8] BWEB[9] BWEB[10] BWEB[11] BWEB[12] BWEB[13] BWEB[14] BWEB[15]
+ BWEB[16] VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD
+ VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD
+ VLO_VXDD VLO_VXDD CKD D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] D[8] D[9] D[10]
+ D[11] D[12] D[13] D[14] D[15] D[16] VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD
+ VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD
+ VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD GBL[0] GBL[1] GBL[2] GBL[3]
+ GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13]
+ GBL[14] GBL[15] GBL[16] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5]
+ GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14]
+ GBLB[15] GBLB[16] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9]
+ GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GWB[0] GWB[1] GWB[2] GWB[3]
+ GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13]
+ GWB[14] GWB[15] GWB[16] SLP_BUF SLP_BUF PDO Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6]
+ Q[7] Q[8] Q[9] Q[10] Q[11] Q[12] Q[13] Q[14] Q[15] Q[16] SLP_Q VXDDHD VDD VSS
+ VLO WLP_SAEB SLP_LBACK VXDDHD VDD VLO_VXDD VXDDHD S1BSVTSWSO8000Y24_MIO_L_DR
XMIO_R AWT2 VLO_VXDD BWEB[19] BWEB[20] BWEB[21] BWEB[22] BWEB[23] BWEB[24]
+ BWEB[25] BWEB[26] BWEB[27] BWEB[28] BWEB[29] BWEB[30] BWEB[31] BWEB[32]
+ BWEB[33] BWEB[34] BWEB[35] VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD
+ VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD
+ VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD CKD D[19] D[20] D[21] D[22] D[23] D[24]
+ D[25] D[26] D[27] D[28] D[29] D[30] D[31] D[32] D[33] D[34] D[35] VLO_VXDD
+ VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD
+ VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBLB[19]
+ GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27]
+ GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GW[19]
+ GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30]
+ GW[31] GW[32] GW[33] GW[34] GW[35] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23]
+ GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32]
+ GWB[33] GWB[34] GWB[35] SLP_BUF SLP_BUF PDO Q[19] Q[20] Q[21] Q[22] Q[23]
+ Q[24] Q[25] Q[26] Q[27] Q[28] Q[29] Q[30] Q[31] Q[32] Q[33] Q[34] Q[35] SLP_Q
+ VXDDHD VDD VSS VLO WLP_SAEB SLP_RBACK VXDDHD VDD VLO_VXDD VXDDHD
+ S1BSVTSWSO8000Y24_MIO_R_DR
XCNT_CORE_IO_M16 VLO_VXDD AWT2 VLO_VXDD VLO_VXDD BLTRKWLDRV CEB VLO_VXDD CKD CLK
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5]
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0]
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] VHI_VXDD
+ VLO_VXDD RE WE TK VLO_VXDD TRKBL VXDDHD VDD VHI VLO VSS WEB VLO_VXDD WLP_SAE
+ WLP_SAEB WLP_SAE_TK VLO_VXDD VLO_VXDD VLO_VXDD A[4] A[5] A[6] A[7] A[8] A[9]
+ A[10] A[11] A[12] A[13] A[14] VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD
+ VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD A[0] A[1] A[2] A[3]
+ YL[0] YL[1] VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD VLO_VXDD DSLP_BUF SD SD_BUF
+ SLP SLP_BUF SLP_LBACK SLP_LCTRL SLP_Q SLP_RBACK BWEB[17] BWEB[18] VLO_VXDD
+ VLO_VXDD D[17] D[18] VLO_VXDD VLO_VXDD GBL[17] GBL[18] GBLB[17] GBLB[18]
+ GW[17] GW[18] GWB[17] GWB[18] Q[17] Q[18] VXDDHD VDD VLO_VXDD VLO_VXDD
+ VHI_VXDD S1BSVTSWSO8000Y24_CNT_CORE_IO_DR
XTOPEDGE VXDDHD VDD VSS WLP_SAE WLP_SAE_TK S1BSVTSWSO8000Y24_TOP_EDGE
XD_WEB WEB VSS S1BSVTSWSO8000Y24_DIO
XD_CEB CEB VSS S1BSVTSWSO8000Y24_DIO
XD_CLK CLK VSS S1BSVTSWSO8000Y24_DIO
XD_SLP SLP VSS S1BSVTSWSO8000Y24_DIO
XD_SD SD VSS S1BSVTSWSO8000Y24_DIO
XD_A0 A[0] VSS S1BSVTSWSO8000Y24_DIO
XD_A1 A[1] VSS S1BSVTSWSO8000Y24_DIO
XD_A2 A[2] VSS S1BSVTSWSO8000Y24_DIO
XD_A3 A[3] VSS S1BSVTSWSO8000Y24_DIO
XD_A4 A[4] VSS S1BSVTSWSO8000Y24_DIO
XD_A5 A[5] VSS S1BSVTSWSO8000Y24_DIO
XD_A6 A[6] VSS S1BSVTSWSO8000Y24_DIO
XD_A7 A[7] VSS S1BSVTSWSO8000Y24_DIO
XD_A8 A[8] VSS S1BSVTSWSO8000Y24_DIO
XD_A9 A[9] VSS S1BSVTSWSO8000Y24_DIO
XD_A10 A[10] VSS S1BSVTSWSO8000Y24_DIO
XD_A11 A[11] VSS S1BSVTSWSO8000Y24_DIO
XD_A12 A[12] VSS S1BSVTSWSO8000Y24_DIO
XD_A13 A[13] VSS S1BSVTSWSO8000Y24_DIO
XD_A14 A[14] VSS S1BSVTSWSO8000Y24_DIO
XD_D0 D[0] VSS S1BSVTSWSO8000Y24_DIO
XD_D1 D[1] VSS S1BSVTSWSO8000Y24_DIO
XD_D2 D[2] VSS S1BSVTSWSO8000Y24_DIO
XD_D3 D[3] VSS S1BSVTSWSO8000Y24_DIO
XD_D4 D[4] VSS S1BSVTSWSO8000Y24_DIO
XD_D5 D[5] VSS S1BSVTSWSO8000Y24_DIO
XD_D6 D[6] VSS S1BSVTSWSO8000Y24_DIO
XD_D7 D[7] VSS S1BSVTSWSO8000Y24_DIO
XD_D8 D[8] VSS S1BSVTSWSO8000Y24_DIO
XD_D9 D[9] VSS S1BSVTSWSO8000Y24_DIO
XD_D10 D[10] VSS S1BSVTSWSO8000Y24_DIO
XD_D11 D[11] VSS S1BSVTSWSO8000Y24_DIO
XD_D12 D[12] VSS S1BSVTSWSO8000Y24_DIO
XD_D13 D[13] VSS S1BSVTSWSO8000Y24_DIO
XD_D14 D[14] VSS S1BSVTSWSO8000Y24_DIO
XD_D15 D[15] VSS S1BSVTSWSO8000Y24_DIO
XD_D16 D[16] VSS S1BSVTSWSO8000Y24_DIO
XD_D17 D[17] VSS S1BSVTSWSO8000Y24_DIO
XD_D18 D[18] VSS S1BSVTSWSO8000Y24_DIO
XD_D19 D[19] VSS S1BSVTSWSO8000Y24_DIO
XD_D20 D[20] VSS S1BSVTSWSO8000Y24_DIO
XD_D21 D[21] VSS S1BSVTSWSO8000Y24_DIO
XD_D22 D[22] VSS S1BSVTSWSO8000Y24_DIO
XD_D23 D[23] VSS S1BSVTSWSO8000Y24_DIO
XD_D24 D[24] VSS S1BSVTSWSO8000Y24_DIO
XD_D25 D[25] VSS S1BSVTSWSO8000Y24_DIO
XD_D26 D[26] VSS S1BSVTSWSO8000Y24_DIO
XD_D27 D[27] VSS S1BSVTSWSO8000Y24_DIO
XD_D28 D[28] VSS S1BSVTSWSO8000Y24_DIO
XD_D29 D[29] VSS S1BSVTSWSO8000Y24_DIO
XD_D30 D[30] VSS S1BSVTSWSO8000Y24_DIO
XD_D31 D[31] VSS S1BSVTSWSO8000Y24_DIO
XD_D32 D[32] VSS S1BSVTSWSO8000Y24_DIO
XD_D33 D[33] VSS S1BSVTSWSO8000Y24_DIO
XD_D34 D[34] VSS S1BSVTSWSO8000Y24_DIO
XD_D35 D[35] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB0 BWEB[0] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB1 BWEB[1] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB2 BWEB[2] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB3 BWEB[3] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB4 BWEB[4] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB5 BWEB[5] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB6 BWEB[6] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB7 BWEB[7] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB8 BWEB[8] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB9 BWEB[9] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB10 BWEB[10] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB11 BWEB[11] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB12 BWEB[12] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB13 BWEB[13] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB14 BWEB[14] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB15 BWEB[15] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB16 BWEB[16] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB17 BWEB[17] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB18 BWEB[18] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB19 BWEB[19] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB20 BWEB[20] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB21 BWEB[21] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB22 BWEB[22] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB23 BWEB[23] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB24 BWEB[24] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB25 BWEB[25] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB26 BWEB[26] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB27 BWEB[27] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB28 BWEB[28] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB29 BWEB[29] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB30 BWEB[30] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB31 BWEB[31] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB32 BWEB[32] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB33 BWEB[33] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB34 BWEB[34] VSS S1BSVTSWSO8000Y24_DIO
XD_BWEB35 BWEB[35] VSS S1BSVTSWSO8000Y24_DIO
.ENDS

